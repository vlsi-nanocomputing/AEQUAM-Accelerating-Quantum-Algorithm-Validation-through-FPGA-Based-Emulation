LIBRARY IEEE;
USE WORK.COMB_ADDER;
USE IEEE.NUMERIC_STD.ALL;

ARCHITECTURE behavioral OF comb_adder IS 

SIGNAL RESULT : STD_LOGIC_VECTOR(K DOWNTO 0);


BEGIN

	RESULT <= STD_LOGIC_VECTOR ( SIGNED(COMB_ADD_IN_A) + SIGNED(COMB_ADD_IN_B) + TO_SIGNED(0,K)&COMB_ADD_IN_CIN);
	
	COMB_ADD_OUT_RES <= RESULT (K DOWNTO 1);

END behavioral;