library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_64_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_64_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_32 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_33 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_34 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_35 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_36 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_37 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_38 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_39 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_40 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_41 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_42 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_43 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_44 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_45 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_46 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_47 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_48 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_49 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_50 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_51 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_52 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_53 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_54 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_55 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_56 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_57 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_58 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_59 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_60 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_61 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_62 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_63 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_SEL : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		MUX_64_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_64_1 IS

BEGIN

	MUX_64_1_OUT_RES <= 
				MUX_64_1_IN_0 WHEN MUX_64_1_IN_SEL = "000000" ELSE
				MUX_64_1_IN_1 WHEN MUX_64_1_IN_SEL = "000001" ELSE
				MUX_64_1_IN_2 WHEN MUX_64_1_IN_SEL = "000010" ELSE
				MUX_64_1_IN_3 WHEN MUX_64_1_IN_SEL = "000011" ELSE
				MUX_64_1_IN_4 WHEN MUX_64_1_IN_SEL = "000100" ELSE
				MUX_64_1_IN_5 WHEN MUX_64_1_IN_SEL = "000101" ELSE
				MUX_64_1_IN_6 WHEN MUX_64_1_IN_SEL = "000110" ELSE
				MUX_64_1_IN_7 WHEN MUX_64_1_IN_SEL = "000111" ELSE
				MUX_64_1_IN_8 WHEN MUX_64_1_IN_SEL = "001000" ELSE
				MUX_64_1_IN_9 WHEN MUX_64_1_IN_SEL = "001001" ELSE
				MUX_64_1_IN_10 WHEN MUX_64_1_IN_SEL = "001010" ELSE
				MUX_64_1_IN_11 WHEN MUX_64_1_IN_SEL = "001011" ELSE
				MUX_64_1_IN_12 WHEN MUX_64_1_IN_SEL = "001100" ELSE
				MUX_64_1_IN_13 WHEN MUX_64_1_IN_SEL = "001101" ELSE
				MUX_64_1_IN_14 WHEN MUX_64_1_IN_SEL = "001110" ELSE
				MUX_64_1_IN_15 WHEN MUX_64_1_IN_SEL = "001111" ELSE
				MUX_64_1_IN_16 WHEN MUX_64_1_IN_SEL = "010000" ELSE
				MUX_64_1_IN_17 WHEN MUX_64_1_IN_SEL = "010001" ELSE
				MUX_64_1_IN_18 WHEN MUX_64_1_IN_SEL = "010010" ELSE
				MUX_64_1_IN_19 WHEN MUX_64_1_IN_SEL = "010011" ELSE
				MUX_64_1_IN_20 WHEN MUX_64_1_IN_SEL = "010100" ELSE
				MUX_64_1_IN_21 WHEN MUX_64_1_IN_SEL = "010101" ELSE
				MUX_64_1_IN_22 WHEN MUX_64_1_IN_SEL = "010110" ELSE
				MUX_64_1_IN_23 WHEN MUX_64_1_IN_SEL = "010111" ELSE
				MUX_64_1_IN_24 WHEN MUX_64_1_IN_SEL = "011000" ELSE
				MUX_64_1_IN_25 WHEN MUX_64_1_IN_SEL = "011001" ELSE
				MUX_64_1_IN_26 WHEN MUX_64_1_IN_SEL = "011010" ELSE
				MUX_64_1_IN_27 WHEN MUX_64_1_IN_SEL = "011011" ELSE
				MUX_64_1_IN_28 WHEN MUX_64_1_IN_SEL = "011100" ELSE
				MUX_64_1_IN_29 WHEN MUX_64_1_IN_SEL = "011101" ELSE
				MUX_64_1_IN_30 WHEN MUX_64_1_IN_SEL = "011110" ELSE
				MUX_64_1_IN_31 WHEN MUX_64_1_IN_SEL = "011111" ELSE
				MUX_64_1_IN_32 WHEN MUX_64_1_IN_SEL = "100000" ELSE
				MUX_64_1_IN_33 WHEN MUX_64_1_IN_SEL = "100001" ELSE
				MUX_64_1_IN_34 WHEN MUX_64_1_IN_SEL = "100010" ELSE
				MUX_64_1_IN_35 WHEN MUX_64_1_IN_SEL = "100011" ELSE
				MUX_64_1_IN_36 WHEN MUX_64_1_IN_SEL = "100100" ELSE
				MUX_64_1_IN_37 WHEN MUX_64_1_IN_SEL = "100101" ELSE
				MUX_64_1_IN_38 WHEN MUX_64_1_IN_SEL = "100110" ELSE
				MUX_64_1_IN_39 WHEN MUX_64_1_IN_SEL = "100111" ELSE
				MUX_64_1_IN_40 WHEN MUX_64_1_IN_SEL = "101000" ELSE
				MUX_64_1_IN_41 WHEN MUX_64_1_IN_SEL = "101001" ELSE
				MUX_64_1_IN_42 WHEN MUX_64_1_IN_SEL = "101010" ELSE
				MUX_64_1_IN_43 WHEN MUX_64_1_IN_SEL = "101011" ELSE
				MUX_64_1_IN_44 WHEN MUX_64_1_IN_SEL = "101100" ELSE
				MUX_64_1_IN_45 WHEN MUX_64_1_IN_SEL = "101101" ELSE
				MUX_64_1_IN_46 WHEN MUX_64_1_IN_SEL = "101110" ELSE
				MUX_64_1_IN_47 WHEN MUX_64_1_IN_SEL = "101111" ELSE
				MUX_64_1_IN_48 WHEN MUX_64_1_IN_SEL = "110000" ELSE
				MUX_64_1_IN_49 WHEN MUX_64_1_IN_SEL = "110001" ELSE
				MUX_64_1_IN_50 WHEN MUX_64_1_IN_SEL = "110010" ELSE
				MUX_64_1_IN_51 WHEN MUX_64_1_IN_SEL = "110011" ELSE
				MUX_64_1_IN_52 WHEN MUX_64_1_IN_SEL = "110100" ELSE
				MUX_64_1_IN_53 WHEN MUX_64_1_IN_SEL = "110101" ELSE
				MUX_64_1_IN_54 WHEN MUX_64_1_IN_SEL = "110110" ELSE
				MUX_64_1_IN_55 WHEN MUX_64_1_IN_SEL = "110111" ELSE
				MUX_64_1_IN_56 WHEN MUX_64_1_IN_SEL = "111000" ELSE
				MUX_64_1_IN_57 WHEN MUX_64_1_IN_SEL = "111001" ELSE
				MUX_64_1_IN_58 WHEN MUX_64_1_IN_SEL = "111010" ELSE
				MUX_64_1_IN_59 WHEN MUX_64_1_IN_SEL = "111011" ELSE
				MUX_64_1_IN_60 WHEN MUX_64_1_IN_SEL = "111100" ELSE
				MUX_64_1_IN_61 WHEN MUX_64_1_IN_SEL = "111101" ELSE
				MUX_64_1_IN_62 WHEN MUX_64_1_IN_SEL = "111110" ELSE
				MUX_64_1_IN_63 WHEN MUX_64_1_IN_SEL = "111111" ELSE
				(OTHERS => '0');


END behavioral;