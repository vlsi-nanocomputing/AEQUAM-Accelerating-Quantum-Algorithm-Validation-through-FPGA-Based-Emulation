LIBRARY IEEE;
USE WORK.MULTIPLIER;
USE IEEE.NUMERIC_STD.ALL;

ARCHITECTURE behavioral OF multiplier IS

BEGIN

	MULTIPLIER_OUT_RES <= STD_LOGIC_VECTOR( SIGNED( MULTIPLIER_IN_A ) * SIGNED( MULTIPLIER_IN_B ) );

END behavioral;