library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY QEP_N_10_W_0_S_0 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		QEP_N_10_W_0_S_0_IN_START : IN STD_LOGIC;
		QEP_N_10_W_0_S_0_IN_QTGT : IN STD_LOGIC_VECTOR (3 DOWNTO 0);  
		QEP_N_10_W_0_S_0_IN_CTRL_MASK : IN STD_LOGIC_VECTOR(1023 DOWNTO 0);
		QEP_N_10_W_0_S_0_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		QEP_N_10_W_0_S_0_IN_SIN : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_10_W_0_S_0_IN_COS : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_10_W_0_S_0_IN_OUT_STATE_SEL : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		QEP_N_10_W_0_S_0_IN_REAL_IMAG_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		QEP_N_10_W_0_S_0_IN_CLK : IN STD_LOGIC;
		QEP_N_10_W_0_S_0_IN_CLEAR : IN STD_LOGIC;
		QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF : IN STD_LOGIC;
		QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE : IN STD_LOGIC;
		QEP_N_10_W_0_S_0_OUT_DONE : OUT STD_LOGIC;
		QEP_N_10_W_0_S_0_OUT_DATA : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;
ARCHITECTURE generated OF QEP_N_10_W_0_S_0 IS
COMPONENT multiplexer_2_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_2_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		MUX_2_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_10_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_10_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_10_1_IN_SEL : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		MUX_10_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_1024_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_1024_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_32 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_33 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_34 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_35 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_36 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_37 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_38 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_39 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_40 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_41 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_42 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_43 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_44 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_45 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_46 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_47 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_48 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_49 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_50 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_51 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_52 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_53 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_54 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_55 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_56 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_57 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_58 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_59 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_60 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_61 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_62 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_63 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_64 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_65 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_66 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_67 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_68 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_69 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_70 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_71 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_72 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_73 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_74 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_75 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_76 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_77 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_78 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_79 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_80 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_81 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_82 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_83 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_84 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_85 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_86 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_87 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_88 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_89 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_90 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_91 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_92 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_93 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_94 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_95 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_96 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_97 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_98 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_99 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_100 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_101 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_102 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_103 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_104 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_105 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_106 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_107 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_108 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_109 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_110 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_111 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_112 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_113 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_114 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_115 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_116 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_117 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_118 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_119 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_120 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_121 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_122 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_123 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_124 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_125 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_126 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_127 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_128 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_129 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_130 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_131 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_132 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_133 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_134 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_135 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_136 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_137 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_138 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_139 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_140 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_141 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_142 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_143 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_144 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_145 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_146 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_147 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_148 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_149 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_150 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_151 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_152 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_153 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_154 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_155 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_156 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_157 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_158 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_159 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_160 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_161 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_162 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_163 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_164 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_165 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_166 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_167 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_168 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_169 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_170 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_171 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_172 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_173 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_174 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_175 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_176 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_177 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_178 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_179 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_180 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_181 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_182 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_183 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_184 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_185 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_186 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_187 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_188 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_189 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_190 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_191 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_192 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_193 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_194 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_195 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_196 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_197 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_198 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_199 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_200 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_201 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_202 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_203 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_204 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_205 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_206 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_207 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_208 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_209 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_210 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_211 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_212 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_213 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_214 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_215 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_216 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_217 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_218 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_219 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_220 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_221 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_222 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_223 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_224 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_225 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_226 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_227 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_228 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_229 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_230 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_231 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_232 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_233 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_234 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_235 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_236 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_237 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_238 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_239 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_240 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_241 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_242 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_243 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_244 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_245 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_246 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_247 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_248 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_249 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_250 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_251 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_252 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_253 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_254 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_255 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_256 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_257 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_258 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_259 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_260 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_261 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_262 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_263 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_264 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_265 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_266 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_267 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_268 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_269 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_270 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_271 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_272 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_273 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_274 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_275 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_276 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_277 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_278 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_279 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_280 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_281 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_282 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_283 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_284 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_285 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_286 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_287 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_288 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_289 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_290 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_291 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_292 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_293 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_294 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_295 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_296 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_297 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_298 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_299 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_300 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_301 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_302 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_303 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_304 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_305 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_306 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_307 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_308 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_309 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_310 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_311 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_312 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_313 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_314 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_315 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_316 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_317 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_318 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_319 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_320 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_321 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_322 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_323 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_324 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_325 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_326 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_327 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_328 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_329 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_330 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_331 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_332 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_333 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_334 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_335 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_336 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_337 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_338 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_339 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_340 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_341 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_342 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_343 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_344 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_345 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_346 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_347 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_348 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_349 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_350 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_351 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_352 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_353 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_354 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_355 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_356 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_357 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_358 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_359 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_360 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_361 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_362 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_363 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_364 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_365 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_366 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_367 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_368 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_369 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_370 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_371 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_372 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_373 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_374 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_375 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_376 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_377 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_378 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_379 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_380 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_381 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_382 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_383 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_384 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_385 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_386 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_387 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_388 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_389 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_390 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_391 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_392 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_393 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_394 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_395 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_396 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_397 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_398 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_399 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_400 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_401 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_402 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_403 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_404 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_405 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_406 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_407 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_408 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_409 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_410 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_411 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_412 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_413 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_414 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_415 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_416 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_417 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_418 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_419 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_420 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_421 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_422 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_423 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_424 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_425 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_426 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_427 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_428 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_429 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_430 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_431 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_432 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_433 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_434 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_435 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_436 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_437 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_438 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_439 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_440 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_441 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_442 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_443 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_444 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_445 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_446 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_447 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_448 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_449 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_450 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_451 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_452 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_453 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_454 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_455 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_456 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_457 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_458 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_459 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_460 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_461 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_462 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_463 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_464 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_465 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_466 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_467 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_468 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_469 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_470 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_471 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_472 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_473 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_474 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_475 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_476 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_477 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_478 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_479 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_480 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_481 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_482 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_483 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_484 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_485 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_486 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_487 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_488 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_489 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_490 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_491 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_492 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_493 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_494 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_495 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_496 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_497 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_498 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_499 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_500 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_501 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_502 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_503 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_504 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_505 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_506 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_507 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_508 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_509 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_510 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_511 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_512 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_513 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_514 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_515 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_516 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_517 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_518 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_519 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_520 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_521 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_522 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_523 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_524 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_525 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_526 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_527 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_528 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_529 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_530 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_531 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_532 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_533 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_534 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_535 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_536 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_537 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_538 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_539 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_540 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_541 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_542 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_543 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_544 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_545 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_546 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_547 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_548 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_549 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_550 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_551 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_552 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_553 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_554 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_555 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_556 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_557 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_558 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_559 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_560 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_561 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_562 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_563 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_564 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_565 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_566 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_567 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_568 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_569 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_570 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_571 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_572 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_573 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_574 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_575 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_576 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_577 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_578 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_579 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_580 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_581 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_582 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_583 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_584 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_585 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_586 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_587 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_588 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_589 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_590 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_591 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_592 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_593 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_594 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_595 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_596 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_597 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_598 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_599 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_600 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_601 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_602 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_603 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_604 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_605 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_606 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_607 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_608 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_609 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_610 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_611 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_612 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_613 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_614 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_615 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_616 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_617 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_618 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_619 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_620 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_621 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_622 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_623 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_624 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_625 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_626 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_627 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_628 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_629 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_630 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_631 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_632 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_633 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_634 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_635 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_636 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_637 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_638 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_639 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_640 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_641 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_642 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_643 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_644 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_645 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_646 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_647 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_648 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_649 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_650 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_651 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_652 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_653 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_654 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_655 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_656 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_657 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_658 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_659 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_660 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_661 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_662 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_663 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_664 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_665 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_666 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_667 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_668 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_669 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_670 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_671 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_672 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_673 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_674 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_675 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_676 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_677 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_678 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_679 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_680 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_681 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_682 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_683 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_684 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_685 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_686 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_687 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_688 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_689 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_690 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_691 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_692 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_693 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_694 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_695 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_696 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_697 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_698 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_699 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_700 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_701 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_702 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_703 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_704 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_705 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_706 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_707 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_708 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_709 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_710 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_711 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_712 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_713 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_714 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_715 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_716 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_717 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_718 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_719 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_720 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_721 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_722 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_723 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_724 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_725 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_726 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_727 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_728 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_729 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_730 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_731 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_732 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_733 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_734 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_735 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_736 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_737 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_738 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_739 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_740 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_741 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_742 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_743 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_744 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_745 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_746 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_747 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_748 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_749 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_750 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_751 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_752 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_753 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_754 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_755 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_756 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_757 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_758 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_759 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_760 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_761 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_762 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_763 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_764 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_765 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_766 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_767 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_768 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_769 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_770 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_771 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_772 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_773 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_774 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_775 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_776 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_777 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_778 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_779 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_780 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_781 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_782 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_783 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_784 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_785 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_786 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_787 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_788 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_789 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_790 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_791 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_792 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_793 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_794 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_795 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_796 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_797 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_798 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_799 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_800 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_801 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_802 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_803 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_804 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_805 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_806 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_807 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_808 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_809 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_810 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_811 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_812 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_813 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_814 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_815 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_816 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_817 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_818 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_819 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_820 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_821 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_822 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_823 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_824 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_825 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_826 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_827 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_828 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_829 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_830 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_831 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_832 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_833 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_834 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_835 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_836 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_837 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_838 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_839 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_840 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_841 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_842 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_843 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_844 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_845 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_846 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_847 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_848 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_849 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_850 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_851 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_852 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_853 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_854 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_855 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_856 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_857 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_858 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_859 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_860 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_861 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_862 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_863 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_864 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_865 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_866 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_867 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_868 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_869 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_870 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_871 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_872 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_873 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_874 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_875 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_876 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_877 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_878 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_879 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_880 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_881 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_882 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_883 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_884 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_885 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_886 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_887 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_888 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_889 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_890 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_891 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_892 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_893 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_894 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_895 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_896 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_897 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_898 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_899 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_900 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_901 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_902 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_903 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_904 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_905 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_906 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_907 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_908 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_909 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_910 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_911 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_912 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_913 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_914 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_915 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_916 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_917 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_918 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_919 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_920 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_921 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_922 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_923 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_924 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_925 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_926 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_927 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_928 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_929 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_930 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_931 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_932 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_933 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_934 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_935 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_936 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_937 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_938 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_939 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_940 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_941 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_942 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_943 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_944 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_945 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_946 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_947 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_948 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_949 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_950 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_951 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_952 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_953 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_954 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_955 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_956 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_957 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_958 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_959 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_960 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_961 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_962 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_963 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_964 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_965 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_966 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_967 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_968 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_969 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_970 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_971 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_972 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_973 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_974 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_975 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_976 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_977 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_978 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_979 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_980 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_981 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_982 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_983 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_984 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_985 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_986 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_987 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_988 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_989 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_990 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_991 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_992 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_993 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_994 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_995 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_996 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_997 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_998 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_999 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1000 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1001 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1002 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1003 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1004 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1005 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1006 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1007 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1008 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1009 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1010 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1011 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1012 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1013 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1014 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1015 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1016 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1017 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1018 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1019 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1020 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1021 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1022 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1023 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_SEL : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		MUX_1024_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register_clear_1 IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT datapath is
    GENERIC (K : INTEGER := 20);	--K represents the chosen parallelism
	PORT(
		--Data signals
		DATAPATH_IN_A : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_B : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_SINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_COSINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_PIPE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_LD : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_MUX_CTRL : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
		DATAPATH_IN_SUB : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		DATAPATH_IN_SAVED : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_CLEAR : IN STD_LOGIC;
		DATAPATH_IN_CLK : IN STD_LOGIC;
		DATAPATH_OUT_A : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_OUT_B : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0));
END COMPONENT;
COMPONENT control_unit IS
 	PORT (
		--Input signals
		CONTROL_UNIT_IN_START : IN STD_LOGIC;
		CONTROL_UNIT_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CONTROL_UNIT_IN_CLK : IN STD_LOGIC;
		CONTROL_UNIT_IN_CLEAR : IN STD_LOGIC;
		CONTROL_UNIT_OUT_PIPE: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_LD : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_MUX_CTRL : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
		CONTROL_UNIT_OUT_SUB : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		CONTROL_UNIT_OUT_SAVED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_DONE : OUT STD_LOGIC);
END COMPONENT;

SIGNAL TO_STATE_REG_0,TO_STATE_REG_1,TO_STATE_REG_2,TO_STATE_REG_3,TO_STATE_REG_4,TO_STATE_REG_5,TO_STATE_REG_6,TO_STATE_REG_7,TO_STATE_REG_8,TO_STATE_REG_9,TO_STATE_REG_10,TO_STATE_REG_11,TO_STATE_REG_12,TO_STATE_REG_13,TO_STATE_REG_14,TO_STATE_REG_15,TO_STATE_REG_16,TO_STATE_REG_17,TO_STATE_REG_18,TO_STATE_REG_19,TO_STATE_REG_20,TO_STATE_REG_21,TO_STATE_REG_22,TO_STATE_REG_23,TO_STATE_REG_24,TO_STATE_REG_25,TO_STATE_REG_26,TO_STATE_REG_27,TO_STATE_REG_28,TO_STATE_REG_29,TO_STATE_REG_30,TO_STATE_REG_31,TO_STATE_REG_32,TO_STATE_REG_33,TO_STATE_REG_34,TO_STATE_REG_35,TO_STATE_REG_36,TO_STATE_REG_37,TO_STATE_REG_38,TO_STATE_REG_39,TO_STATE_REG_40,TO_STATE_REG_41,TO_STATE_REG_42,TO_STATE_REG_43,TO_STATE_REG_44,TO_STATE_REG_45,TO_STATE_REG_46,TO_STATE_REG_47,TO_STATE_REG_48,TO_STATE_REG_49,TO_STATE_REG_50,TO_STATE_REG_51,TO_STATE_REG_52,TO_STATE_REG_53,TO_STATE_REG_54,TO_STATE_REG_55,TO_STATE_REG_56,TO_STATE_REG_57,TO_STATE_REG_58,TO_STATE_REG_59,TO_STATE_REG_60,TO_STATE_REG_61,TO_STATE_REG_62,TO_STATE_REG_63,TO_STATE_REG_64,TO_STATE_REG_65,TO_STATE_REG_66,TO_STATE_REG_67,TO_STATE_REG_68,TO_STATE_REG_69,TO_STATE_REG_70,TO_STATE_REG_71,TO_STATE_REG_72,TO_STATE_REG_73,TO_STATE_REG_74,TO_STATE_REG_75,TO_STATE_REG_76,TO_STATE_REG_77,TO_STATE_REG_78,TO_STATE_REG_79,TO_STATE_REG_80,TO_STATE_REG_81,TO_STATE_REG_82,TO_STATE_REG_83,TO_STATE_REG_84,TO_STATE_REG_85,TO_STATE_REG_86,TO_STATE_REG_87,TO_STATE_REG_88,TO_STATE_REG_89,TO_STATE_REG_90,TO_STATE_REG_91,TO_STATE_REG_92,TO_STATE_REG_93,TO_STATE_REG_94,TO_STATE_REG_95,TO_STATE_REG_96,TO_STATE_REG_97,TO_STATE_REG_98,TO_STATE_REG_99,TO_STATE_REG_100,TO_STATE_REG_101,TO_STATE_REG_102,TO_STATE_REG_103,TO_STATE_REG_104,TO_STATE_REG_105,TO_STATE_REG_106,TO_STATE_REG_107,TO_STATE_REG_108,TO_STATE_REG_109,TO_STATE_REG_110,TO_STATE_REG_111,TO_STATE_REG_112,TO_STATE_REG_113,TO_STATE_REG_114,TO_STATE_REG_115,TO_STATE_REG_116,TO_STATE_REG_117,TO_STATE_REG_118,TO_STATE_REG_119,TO_STATE_REG_120,TO_STATE_REG_121,TO_STATE_REG_122,TO_STATE_REG_123,TO_STATE_REG_124,TO_STATE_REG_125,TO_STATE_REG_126,TO_STATE_REG_127,TO_STATE_REG_128,TO_STATE_REG_129,TO_STATE_REG_130,TO_STATE_REG_131,TO_STATE_REG_132,TO_STATE_REG_133,TO_STATE_REG_134,TO_STATE_REG_135,TO_STATE_REG_136,TO_STATE_REG_137,TO_STATE_REG_138,TO_STATE_REG_139,TO_STATE_REG_140,TO_STATE_REG_141,TO_STATE_REG_142,TO_STATE_REG_143,TO_STATE_REG_144,TO_STATE_REG_145,TO_STATE_REG_146,TO_STATE_REG_147,TO_STATE_REG_148,TO_STATE_REG_149,TO_STATE_REG_150,TO_STATE_REG_151,TO_STATE_REG_152,TO_STATE_REG_153,TO_STATE_REG_154,TO_STATE_REG_155,TO_STATE_REG_156,TO_STATE_REG_157,TO_STATE_REG_158,TO_STATE_REG_159,TO_STATE_REG_160,TO_STATE_REG_161,TO_STATE_REG_162,TO_STATE_REG_163,TO_STATE_REG_164,TO_STATE_REG_165,TO_STATE_REG_166,TO_STATE_REG_167,TO_STATE_REG_168,TO_STATE_REG_169,TO_STATE_REG_170,TO_STATE_REG_171,TO_STATE_REG_172,TO_STATE_REG_173,TO_STATE_REG_174,TO_STATE_REG_175,TO_STATE_REG_176,TO_STATE_REG_177,TO_STATE_REG_178,TO_STATE_REG_179,TO_STATE_REG_180,TO_STATE_REG_181,TO_STATE_REG_182,TO_STATE_REG_183,TO_STATE_REG_184,TO_STATE_REG_185,TO_STATE_REG_186,TO_STATE_REG_187,TO_STATE_REG_188,TO_STATE_REG_189,TO_STATE_REG_190,TO_STATE_REG_191,TO_STATE_REG_192,TO_STATE_REG_193,TO_STATE_REG_194,TO_STATE_REG_195,TO_STATE_REG_196,TO_STATE_REG_197,TO_STATE_REG_198,TO_STATE_REG_199,TO_STATE_REG_200,TO_STATE_REG_201,TO_STATE_REG_202,TO_STATE_REG_203,TO_STATE_REG_204,TO_STATE_REG_205,TO_STATE_REG_206,TO_STATE_REG_207,TO_STATE_REG_208,TO_STATE_REG_209,TO_STATE_REG_210,TO_STATE_REG_211,TO_STATE_REG_212,TO_STATE_REG_213,TO_STATE_REG_214,TO_STATE_REG_215,TO_STATE_REG_216,TO_STATE_REG_217,TO_STATE_REG_218,TO_STATE_REG_219,TO_STATE_REG_220,TO_STATE_REG_221,TO_STATE_REG_222,TO_STATE_REG_223,TO_STATE_REG_224,TO_STATE_REG_225,TO_STATE_REG_226,TO_STATE_REG_227,TO_STATE_REG_228,TO_STATE_REG_229,TO_STATE_REG_230,TO_STATE_REG_231,TO_STATE_REG_232,TO_STATE_REG_233,TO_STATE_REG_234,TO_STATE_REG_235,TO_STATE_REG_236,TO_STATE_REG_237,TO_STATE_REG_238,TO_STATE_REG_239,TO_STATE_REG_240,TO_STATE_REG_241,TO_STATE_REG_242,TO_STATE_REG_243,TO_STATE_REG_244,TO_STATE_REG_245,TO_STATE_REG_246,TO_STATE_REG_247,TO_STATE_REG_248,TO_STATE_REG_249,TO_STATE_REG_250,TO_STATE_REG_251,TO_STATE_REG_252,TO_STATE_REG_253,TO_STATE_REG_254,TO_STATE_REG_255,TO_STATE_REG_256,TO_STATE_REG_257,TO_STATE_REG_258,TO_STATE_REG_259,TO_STATE_REG_260,TO_STATE_REG_261,TO_STATE_REG_262,TO_STATE_REG_263,TO_STATE_REG_264,TO_STATE_REG_265,TO_STATE_REG_266,TO_STATE_REG_267,TO_STATE_REG_268,TO_STATE_REG_269,TO_STATE_REG_270,TO_STATE_REG_271,TO_STATE_REG_272,TO_STATE_REG_273,TO_STATE_REG_274,TO_STATE_REG_275,TO_STATE_REG_276,TO_STATE_REG_277,TO_STATE_REG_278,TO_STATE_REG_279,TO_STATE_REG_280,TO_STATE_REG_281,TO_STATE_REG_282,TO_STATE_REG_283,TO_STATE_REG_284,TO_STATE_REG_285,TO_STATE_REG_286,TO_STATE_REG_287,TO_STATE_REG_288,TO_STATE_REG_289,TO_STATE_REG_290,TO_STATE_REG_291,TO_STATE_REG_292,TO_STATE_REG_293,TO_STATE_REG_294,TO_STATE_REG_295,TO_STATE_REG_296,TO_STATE_REG_297,TO_STATE_REG_298,TO_STATE_REG_299,TO_STATE_REG_300,TO_STATE_REG_301,TO_STATE_REG_302,TO_STATE_REG_303,TO_STATE_REG_304,TO_STATE_REG_305,TO_STATE_REG_306,TO_STATE_REG_307,TO_STATE_REG_308,TO_STATE_REG_309,TO_STATE_REG_310,TO_STATE_REG_311,TO_STATE_REG_312,TO_STATE_REG_313,TO_STATE_REG_314,TO_STATE_REG_315,TO_STATE_REG_316,TO_STATE_REG_317,TO_STATE_REG_318,TO_STATE_REG_319,TO_STATE_REG_320,TO_STATE_REG_321,TO_STATE_REG_322,TO_STATE_REG_323,TO_STATE_REG_324,TO_STATE_REG_325,TO_STATE_REG_326,TO_STATE_REG_327,TO_STATE_REG_328,TO_STATE_REG_329,TO_STATE_REG_330,TO_STATE_REG_331,TO_STATE_REG_332,TO_STATE_REG_333,TO_STATE_REG_334,TO_STATE_REG_335,TO_STATE_REG_336,TO_STATE_REG_337,TO_STATE_REG_338,TO_STATE_REG_339,TO_STATE_REG_340,TO_STATE_REG_341,TO_STATE_REG_342,TO_STATE_REG_343,TO_STATE_REG_344,TO_STATE_REG_345,TO_STATE_REG_346,TO_STATE_REG_347,TO_STATE_REG_348,TO_STATE_REG_349,TO_STATE_REG_350,TO_STATE_REG_351,TO_STATE_REG_352,TO_STATE_REG_353,TO_STATE_REG_354,TO_STATE_REG_355,TO_STATE_REG_356,TO_STATE_REG_357,TO_STATE_REG_358,TO_STATE_REG_359,TO_STATE_REG_360,TO_STATE_REG_361,TO_STATE_REG_362,TO_STATE_REG_363,TO_STATE_REG_364,TO_STATE_REG_365,TO_STATE_REG_366,TO_STATE_REG_367,TO_STATE_REG_368,TO_STATE_REG_369,TO_STATE_REG_370,TO_STATE_REG_371,TO_STATE_REG_372,TO_STATE_REG_373,TO_STATE_REG_374,TO_STATE_REG_375,TO_STATE_REG_376,TO_STATE_REG_377,TO_STATE_REG_378,TO_STATE_REG_379,TO_STATE_REG_380,TO_STATE_REG_381,TO_STATE_REG_382,TO_STATE_REG_383,TO_STATE_REG_384,TO_STATE_REG_385,TO_STATE_REG_386,TO_STATE_REG_387,TO_STATE_REG_388,TO_STATE_REG_389,TO_STATE_REG_390,TO_STATE_REG_391,TO_STATE_REG_392,TO_STATE_REG_393,TO_STATE_REG_394,TO_STATE_REG_395,TO_STATE_REG_396,TO_STATE_REG_397,TO_STATE_REG_398,TO_STATE_REG_399,TO_STATE_REG_400,TO_STATE_REG_401,TO_STATE_REG_402,TO_STATE_REG_403,TO_STATE_REG_404,TO_STATE_REG_405,TO_STATE_REG_406,TO_STATE_REG_407,TO_STATE_REG_408,TO_STATE_REG_409,TO_STATE_REG_410,TO_STATE_REG_411,TO_STATE_REG_412,TO_STATE_REG_413,TO_STATE_REG_414,TO_STATE_REG_415,TO_STATE_REG_416,TO_STATE_REG_417,TO_STATE_REG_418,TO_STATE_REG_419,TO_STATE_REG_420,TO_STATE_REG_421,TO_STATE_REG_422,TO_STATE_REG_423,TO_STATE_REG_424,TO_STATE_REG_425,TO_STATE_REG_426,TO_STATE_REG_427,TO_STATE_REG_428,TO_STATE_REG_429,TO_STATE_REG_430,TO_STATE_REG_431,TO_STATE_REG_432,TO_STATE_REG_433,TO_STATE_REG_434,TO_STATE_REG_435,TO_STATE_REG_436,TO_STATE_REG_437,TO_STATE_REG_438,TO_STATE_REG_439,TO_STATE_REG_440,TO_STATE_REG_441,TO_STATE_REG_442,TO_STATE_REG_443,TO_STATE_REG_444,TO_STATE_REG_445,TO_STATE_REG_446,TO_STATE_REG_447,TO_STATE_REG_448,TO_STATE_REG_449,TO_STATE_REG_450,TO_STATE_REG_451,TO_STATE_REG_452,TO_STATE_REG_453,TO_STATE_REG_454,TO_STATE_REG_455,TO_STATE_REG_456,TO_STATE_REG_457,TO_STATE_REG_458,TO_STATE_REG_459,TO_STATE_REG_460,TO_STATE_REG_461,TO_STATE_REG_462,TO_STATE_REG_463,TO_STATE_REG_464,TO_STATE_REG_465,TO_STATE_REG_466,TO_STATE_REG_467,TO_STATE_REG_468,TO_STATE_REG_469,TO_STATE_REG_470,TO_STATE_REG_471,TO_STATE_REG_472,TO_STATE_REG_473,TO_STATE_REG_474,TO_STATE_REG_475,TO_STATE_REG_476,TO_STATE_REG_477,TO_STATE_REG_478,TO_STATE_REG_479,TO_STATE_REG_480,TO_STATE_REG_481,TO_STATE_REG_482,TO_STATE_REG_483,TO_STATE_REG_484,TO_STATE_REG_485,TO_STATE_REG_486,TO_STATE_REG_487,TO_STATE_REG_488,TO_STATE_REG_489,TO_STATE_REG_490,TO_STATE_REG_491,TO_STATE_REG_492,TO_STATE_REG_493,TO_STATE_REG_494,TO_STATE_REG_495,TO_STATE_REG_496,TO_STATE_REG_497,TO_STATE_REG_498,TO_STATE_REG_499,TO_STATE_REG_500,TO_STATE_REG_501,TO_STATE_REG_502,TO_STATE_REG_503,TO_STATE_REG_504,TO_STATE_REG_505,TO_STATE_REG_506,TO_STATE_REG_507,TO_STATE_REG_508,TO_STATE_REG_509,TO_STATE_REG_510,TO_STATE_REG_511,TO_STATE_REG_512,TO_STATE_REG_513,TO_STATE_REG_514,TO_STATE_REG_515,TO_STATE_REG_516,TO_STATE_REG_517,TO_STATE_REG_518,TO_STATE_REG_519,TO_STATE_REG_520,TO_STATE_REG_521,TO_STATE_REG_522,TO_STATE_REG_523,TO_STATE_REG_524,TO_STATE_REG_525,TO_STATE_REG_526,TO_STATE_REG_527,TO_STATE_REG_528,TO_STATE_REG_529,TO_STATE_REG_530,TO_STATE_REG_531,TO_STATE_REG_532,TO_STATE_REG_533,TO_STATE_REG_534,TO_STATE_REG_535,TO_STATE_REG_536,TO_STATE_REG_537,TO_STATE_REG_538,TO_STATE_REG_539,TO_STATE_REG_540,TO_STATE_REG_541,TO_STATE_REG_542,TO_STATE_REG_543,TO_STATE_REG_544,TO_STATE_REG_545,TO_STATE_REG_546,TO_STATE_REG_547,TO_STATE_REG_548,TO_STATE_REG_549,TO_STATE_REG_550,TO_STATE_REG_551,TO_STATE_REG_552,TO_STATE_REG_553,TO_STATE_REG_554,TO_STATE_REG_555,TO_STATE_REG_556,TO_STATE_REG_557,TO_STATE_REG_558,TO_STATE_REG_559,TO_STATE_REG_560,TO_STATE_REG_561,TO_STATE_REG_562,TO_STATE_REG_563,TO_STATE_REG_564,TO_STATE_REG_565,TO_STATE_REG_566,TO_STATE_REG_567,TO_STATE_REG_568,TO_STATE_REG_569,TO_STATE_REG_570,TO_STATE_REG_571,TO_STATE_REG_572,TO_STATE_REG_573,TO_STATE_REG_574,TO_STATE_REG_575,TO_STATE_REG_576,TO_STATE_REG_577,TO_STATE_REG_578,TO_STATE_REG_579,TO_STATE_REG_580,TO_STATE_REG_581,TO_STATE_REG_582,TO_STATE_REG_583,TO_STATE_REG_584,TO_STATE_REG_585,TO_STATE_REG_586,TO_STATE_REG_587,TO_STATE_REG_588,TO_STATE_REG_589,TO_STATE_REG_590,TO_STATE_REG_591,TO_STATE_REG_592,TO_STATE_REG_593,TO_STATE_REG_594,TO_STATE_REG_595,TO_STATE_REG_596,TO_STATE_REG_597,TO_STATE_REG_598,TO_STATE_REG_599,TO_STATE_REG_600,TO_STATE_REG_601,TO_STATE_REG_602,TO_STATE_REG_603,TO_STATE_REG_604,TO_STATE_REG_605,TO_STATE_REG_606,TO_STATE_REG_607,TO_STATE_REG_608,TO_STATE_REG_609,TO_STATE_REG_610,TO_STATE_REG_611,TO_STATE_REG_612,TO_STATE_REG_613,TO_STATE_REG_614,TO_STATE_REG_615,TO_STATE_REG_616,TO_STATE_REG_617,TO_STATE_REG_618,TO_STATE_REG_619,TO_STATE_REG_620,TO_STATE_REG_621,TO_STATE_REG_622,TO_STATE_REG_623,TO_STATE_REG_624,TO_STATE_REG_625,TO_STATE_REG_626,TO_STATE_REG_627,TO_STATE_REG_628,TO_STATE_REG_629,TO_STATE_REG_630,TO_STATE_REG_631,TO_STATE_REG_632,TO_STATE_REG_633,TO_STATE_REG_634,TO_STATE_REG_635,TO_STATE_REG_636,TO_STATE_REG_637,TO_STATE_REG_638,TO_STATE_REG_639,TO_STATE_REG_640,TO_STATE_REG_641,TO_STATE_REG_642,TO_STATE_REG_643,TO_STATE_REG_644,TO_STATE_REG_645,TO_STATE_REG_646,TO_STATE_REG_647,TO_STATE_REG_648,TO_STATE_REG_649,TO_STATE_REG_650,TO_STATE_REG_651,TO_STATE_REG_652,TO_STATE_REG_653,TO_STATE_REG_654,TO_STATE_REG_655,TO_STATE_REG_656,TO_STATE_REG_657,TO_STATE_REG_658,TO_STATE_REG_659,TO_STATE_REG_660,TO_STATE_REG_661,TO_STATE_REG_662,TO_STATE_REG_663,TO_STATE_REG_664,TO_STATE_REG_665,TO_STATE_REG_666,TO_STATE_REG_667,TO_STATE_REG_668,TO_STATE_REG_669,TO_STATE_REG_670,TO_STATE_REG_671,TO_STATE_REG_672,TO_STATE_REG_673,TO_STATE_REG_674,TO_STATE_REG_675,TO_STATE_REG_676,TO_STATE_REG_677,TO_STATE_REG_678,TO_STATE_REG_679,TO_STATE_REG_680,TO_STATE_REG_681,TO_STATE_REG_682,TO_STATE_REG_683,TO_STATE_REG_684,TO_STATE_REG_685,TO_STATE_REG_686,TO_STATE_REG_687,TO_STATE_REG_688,TO_STATE_REG_689,TO_STATE_REG_690,TO_STATE_REG_691,TO_STATE_REG_692,TO_STATE_REG_693,TO_STATE_REG_694,TO_STATE_REG_695,TO_STATE_REG_696,TO_STATE_REG_697,TO_STATE_REG_698,TO_STATE_REG_699,TO_STATE_REG_700,TO_STATE_REG_701,TO_STATE_REG_702,TO_STATE_REG_703,TO_STATE_REG_704,TO_STATE_REG_705,TO_STATE_REG_706,TO_STATE_REG_707,TO_STATE_REG_708,TO_STATE_REG_709,TO_STATE_REG_710,TO_STATE_REG_711,TO_STATE_REG_712,TO_STATE_REG_713,TO_STATE_REG_714,TO_STATE_REG_715,TO_STATE_REG_716,TO_STATE_REG_717,TO_STATE_REG_718,TO_STATE_REG_719,TO_STATE_REG_720,TO_STATE_REG_721,TO_STATE_REG_722,TO_STATE_REG_723,TO_STATE_REG_724,TO_STATE_REG_725,TO_STATE_REG_726,TO_STATE_REG_727,TO_STATE_REG_728,TO_STATE_REG_729,TO_STATE_REG_730,TO_STATE_REG_731,TO_STATE_REG_732,TO_STATE_REG_733,TO_STATE_REG_734,TO_STATE_REG_735,TO_STATE_REG_736,TO_STATE_REG_737,TO_STATE_REG_738,TO_STATE_REG_739,TO_STATE_REG_740,TO_STATE_REG_741,TO_STATE_REG_742,TO_STATE_REG_743,TO_STATE_REG_744,TO_STATE_REG_745,TO_STATE_REG_746,TO_STATE_REG_747,TO_STATE_REG_748,TO_STATE_REG_749,TO_STATE_REG_750,TO_STATE_REG_751,TO_STATE_REG_752,TO_STATE_REG_753,TO_STATE_REG_754,TO_STATE_REG_755,TO_STATE_REG_756,TO_STATE_REG_757,TO_STATE_REG_758,TO_STATE_REG_759,TO_STATE_REG_760,TO_STATE_REG_761,TO_STATE_REG_762,TO_STATE_REG_763,TO_STATE_REG_764,TO_STATE_REG_765,TO_STATE_REG_766,TO_STATE_REG_767,TO_STATE_REG_768,TO_STATE_REG_769,TO_STATE_REG_770,TO_STATE_REG_771,TO_STATE_REG_772,TO_STATE_REG_773,TO_STATE_REG_774,TO_STATE_REG_775,TO_STATE_REG_776,TO_STATE_REG_777,TO_STATE_REG_778,TO_STATE_REG_779,TO_STATE_REG_780,TO_STATE_REG_781,TO_STATE_REG_782,TO_STATE_REG_783,TO_STATE_REG_784,TO_STATE_REG_785,TO_STATE_REG_786,TO_STATE_REG_787,TO_STATE_REG_788,TO_STATE_REG_789,TO_STATE_REG_790,TO_STATE_REG_791,TO_STATE_REG_792,TO_STATE_REG_793,TO_STATE_REG_794,TO_STATE_REG_795,TO_STATE_REG_796,TO_STATE_REG_797,TO_STATE_REG_798,TO_STATE_REG_799,TO_STATE_REG_800,TO_STATE_REG_801,TO_STATE_REG_802,TO_STATE_REG_803,TO_STATE_REG_804,TO_STATE_REG_805,TO_STATE_REG_806,TO_STATE_REG_807,TO_STATE_REG_808,TO_STATE_REG_809,TO_STATE_REG_810,TO_STATE_REG_811,TO_STATE_REG_812,TO_STATE_REG_813,TO_STATE_REG_814,TO_STATE_REG_815,TO_STATE_REG_816,TO_STATE_REG_817,TO_STATE_REG_818,TO_STATE_REG_819,TO_STATE_REG_820,TO_STATE_REG_821,TO_STATE_REG_822,TO_STATE_REG_823,TO_STATE_REG_824,TO_STATE_REG_825,TO_STATE_REG_826,TO_STATE_REG_827,TO_STATE_REG_828,TO_STATE_REG_829,TO_STATE_REG_830,TO_STATE_REG_831,TO_STATE_REG_832,TO_STATE_REG_833,TO_STATE_REG_834,TO_STATE_REG_835,TO_STATE_REG_836,TO_STATE_REG_837,TO_STATE_REG_838,TO_STATE_REG_839,TO_STATE_REG_840,TO_STATE_REG_841,TO_STATE_REG_842,TO_STATE_REG_843,TO_STATE_REG_844,TO_STATE_REG_845,TO_STATE_REG_846,TO_STATE_REG_847,TO_STATE_REG_848,TO_STATE_REG_849,TO_STATE_REG_850,TO_STATE_REG_851,TO_STATE_REG_852,TO_STATE_REG_853,TO_STATE_REG_854,TO_STATE_REG_855,TO_STATE_REG_856,TO_STATE_REG_857,TO_STATE_REG_858,TO_STATE_REG_859,TO_STATE_REG_860,TO_STATE_REG_861,TO_STATE_REG_862,TO_STATE_REG_863,TO_STATE_REG_864,TO_STATE_REG_865,TO_STATE_REG_866,TO_STATE_REG_867,TO_STATE_REG_868,TO_STATE_REG_869,TO_STATE_REG_870,TO_STATE_REG_871,TO_STATE_REG_872,TO_STATE_REG_873,TO_STATE_REG_874,TO_STATE_REG_875,TO_STATE_REG_876,TO_STATE_REG_877,TO_STATE_REG_878,TO_STATE_REG_879,TO_STATE_REG_880,TO_STATE_REG_881,TO_STATE_REG_882,TO_STATE_REG_883,TO_STATE_REG_884,TO_STATE_REG_885,TO_STATE_REG_886,TO_STATE_REG_887,TO_STATE_REG_888,TO_STATE_REG_889,TO_STATE_REG_890,TO_STATE_REG_891,TO_STATE_REG_892,TO_STATE_REG_893,TO_STATE_REG_894,TO_STATE_REG_895,TO_STATE_REG_896,TO_STATE_REG_897,TO_STATE_REG_898,TO_STATE_REG_899,TO_STATE_REG_900,TO_STATE_REG_901,TO_STATE_REG_902,TO_STATE_REG_903,TO_STATE_REG_904,TO_STATE_REG_905,TO_STATE_REG_906,TO_STATE_REG_907,TO_STATE_REG_908,TO_STATE_REG_909,TO_STATE_REG_910,TO_STATE_REG_911,TO_STATE_REG_912,TO_STATE_REG_913,TO_STATE_REG_914,TO_STATE_REG_915,TO_STATE_REG_916,TO_STATE_REG_917,TO_STATE_REG_918,TO_STATE_REG_919,TO_STATE_REG_920,TO_STATE_REG_921,TO_STATE_REG_922,TO_STATE_REG_923,TO_STATE_REG_924,TO_STATE_REG_925,TO_STATE_REG_926,TO_STATE_REG_927,TO_STATE_REG_928,TO_STATE_REG_929,TO_STATE_REG_930,TO_STATE_REG_931,TO_STATE_REG_932,TO_STATE_REG_933,TO_STATE_REG_934,TO_STATE_REG_935,TO_STATE_REG_936,TO_STATE_REG_937,TO_STATE_REG_938,TO_STATE_REG_939,TO_STATE_REG_940,TO_STATE_REG_941,TO_STATE_REG_942,TO_STATE_REG_943,TO_STATE_REG_944,TO_STATE_REG_945,TO_STATE_REG_946,TO_STATE_REG_947,TO_STATE_REG_948,TO_STATE_REG_949,TO_STATE_REG_950,TO_STATE_REG_951,TO_STATE_REG_952,TO_STATE_REG_953,TO_STATE_REG_954,TO_STATE_REG_955,TO_STATE_REG_956,TO_STATE_REG_957,TO_STATE_REG_958,TO_STATE_REG_959,TO_STATE_REG_960,TO_STATE_REG_961,TO_STATE_REG_962,TO_STATE_REG_963,TO_STATE_REG_964,TO_STATE_REG_965,TO_STATE_REG_966,TO_STATE_REG_967,TO_STATE_REG_968,TO_STATE_REG_969,TO_STATE_REG_970,TO_STATE_REG_971,TO_STATE_REG_972,TO_STATE_REG_973,TO_STATE_REG_974,TO_STATE_REG_975,TO_STATE_REG_976,TO_STATE_REG_977,TO_STATE_REG_978,TO_STATE_REG_979,TO_STATE_REG_980,TO_STATE_REG_981,TO_STATE_REG_982,TO_STATE_REG_983,TO_STATE_REG_984,TO_STATE_REG_985,TO_STATE_REG_986,TO_STATE_REG_987,TO_STATE_REG_988,TO_STATE_REG_989,TO_STATE_REG_990,TO_STATE_REG_991,TO_STATE_REG_992,TO_STATE_REG_993,TO_STATE_REG_994,TO_STATE_REG_995,TO_STATE_REG_996,TO_STATE_REG_997,TO_STATE_REG_998,TO_STATE_REG_999,TO_STATE_REG_1000,TO_STATE_REG_1001,TO_STATE_REG_1002,TO_STATE_REG_1003,TO_STATE_REG_1004,TO_STATE_REG_1005,TO_STATE_REG_1006,TO_STATE_REG_1007,TO_STATE_REG_1008,TO_STATE_REG_1009,TO_STATE_REG_1010,TO_STATE_REG_1011,TO_STATE_REG_1012,TO_STATE_REG_1013,TO_STATE_REG_1014,TO_STATE_REG_1015,TO_STATE_REG_1016,TO_STATE_REG_1017,TO_STATE_REG_1018,TO_STATE_REG_1019,TO_STATE_REG_1020,TO_STATE_REG_1021,TO_STATE_REG_1022,TO_STATE_REG_1023: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_STATE_REG_0,FROM_STATE_REG_1,FROM_STATE_REG_2,FROM_STATE_REG_3,FROM_STATE_REG_4,FROM_STATE_REG_5,FROM_STATE_REG_6,FROM_STATE_REG_7,FROM_STATE_REG_8,FROM_STATE_REG_9,FROM_STATE_REG_10,FROM_STATE_REG_11,FROM_STATE_REG_12,FROM_STATE_REG_13,FROM_STATE_REG_14,FROM_STATE_REG_15,FROM_STATE_REG_16,FROM_STATE_REG_17,FROM_STATE_REG_18,FROM_STATE_REG_19,FROM_STATE_REG_20,FROM_STATE_REG_21,FROM_STATE_REG_22,FROM_STATE_REG_23,FROM_STATE_REG_24,FROM_STATE_REG_25,FROM_STATE_REG_26,FROM_STATE_REG_27,FROM_STATE_REG_28,FROM_STATE_REG_29,FROM_STATE_REG_30,FROM_STATE_REG_31,FROM_STATE_REG_32,FROM_STATE_REG_33,FROM_STATE_REG_34,FROM_STATE_REG_35,FROM_STATE_REG_36,FROM_STATE_REG_37,FROM_STATE_REG_38,FROM_STATE_REG_39,FROM_STATE_REG_40,FROM_STATE_REG_41,FROM_STATE_REG_42,FROM_STATE_REG_43,FROM_STATE_REG_44,FROM_STATE_REG_45,FROM_STATE_REG_46,FROM_STATE_REG_47,FROM_STATE_REG_48,FROM_STATE_REG_49,FROM_STATE_REG_50,FROM_STATE_REG_51,FROM_STATE_REG_52,FROM_STATE_REG_53,FROM_STATE_REG_54,FROM_STATE_REG_55,FROM_STATE_REG_56,FROM_STATE_REG_57,FROM_STATE_REG_58,FROM_STATE_REG_59,FROM_STATE_REG_60,FROM_STATE_REG_61,FROM_STATE_REG_62,FROM_STATE_REG_63,FROM_STATE_REG_64,FROM_STATE_REG_65,FROM_STATE_REG_66,FROM_STATE_REG_67,FROM_STATE_REG_68,FROM_STATE_REG_69,FROM_STATE_REG_70,FROM_STATE_REG_71,FROM_STATE_REG_72,FROM_STATE_REG_73,FROM_STATE_REG_74,FROM_STATE_REG_75,FROM_STATE_REG_76,FROM_STATE_REG_77,FROM_STATE_REG_78,FROM_STATE_REG_79,FROM_STATE_REG_80,FROM_STATE_REG_81,FROM_STATE_REG_82,FROM_STATE_REG_83,FROM_STATE_REG_84,FROM_STATE_REG_85,FROM_STATE_REG_86,FROM_STATE_REG_87,FROM_STATE_REG_88,FROM_STATE_REG_89,FROM_STATE_REG_90,FROM_STATE_REG_91,FROM_STATE_REG_92,FROM_STATE_REG_93,FROM_STATE_REG_94,FROM_STATE_REG_95,FROM_STATE_REG_96,FROM_STATE_REG_97,FROM_STATE_REG_98,FROM_STATE_REG_99,FROM_STATE_REG_100,FROM_STATE_REG_101,FROM_STATE_REG_102,FROM_STATE_REG_103,FROM_STATE_REG_104,FROM_STATE_REG_105,FROM_STATE_REG_106,FROM_STATE_REG_107,FROM_STATE_REG_108,FROM_STATE_REG_109,FROM_STATE_REG_110,FROM_STATE_REG_111,FROM_STATE_REG_112,FROM_STATE_REG_113,FROM_STATE_REG_114,FROM_STATE_REG_115,FROM_STATE_REG_116,FROM_STATE_REG_117,FROM_STATE_REG_118,FROM_STATE_REG_119,FROM_STATE_REG_120,FROM_STATE_REG_121,FROM_STATE_REG_122,FROM_STATE_REG_123,FROM_STATE_REG_124,FROM_STATE_REG_125,FROM_STATE_REG_126,FROM_STATE_REG_127,FROM_STATE_REG_128,FROM_STATE_REG_129,FROM_STATE_REG_130,FROM_STATE_REG_131,FROM_STATE_REG_132,FROM_STATE_REG_133,FROM_STATE_REG_134,FROM_STATE_REG_135,FROM_STATE_REG_136,FROM_STATE_REG_137,FROM_STATE_REG_138,FROM_STATE_REG_139,FROM_STATE_REG_140,FROM_STATE_REG_141,FROM_STATE_REG_142,FROM_STATE_REG_143,FROM_STATE_REG_144,FROM_STATE_REG_145,FROM_STATE_REG_146,FROM_STATE_REG_147,FROM_STATE_REG_148,FROM_STATE_REG_149,FROM_STATE_REG_150,FROM_STATE_REG_151,FROM_STATE_REG_152,FROM_STATE_REG_153,FROM_STATE_REG_154,FROM_STATE_REG_155,FROM_STATE_REG_156,FROM_STATE_REG_157,FROM_STATE_REG_158,FROM_STATE_REG_159,FROM_STATE_REG_160,FROM_STATE_REG_161,FROM_STATE_REG_162,FROM_STATE_REG_163,FROM_STATE_REG_164,FROM_STATE_REG_165,FROM_STATE_REG_166,FROM_STATE_REG_167,FROM_STATE_REG_168,FROM_STATE_REG_169,FROM_STATE_REG_170,FROM_STATE_REG_171,FROM_STATE_REG_172,FROM_STATE_REG_173,FROM_STATE_REG_174,FROM_STATE_REG_175,FROM_STATE_REG_176,FROM_STATE_REG_177,FROM_STATE_REG_178,FROM_STATE_REG_179,FROM_STATE_REG_180,FROM_STATE_REG_181,FROM_STATE_REG_182,FROM_STATE_REG_183,FROM_STATE_REG_184,FROM_STATE_REG_185,FROM_STATE_REG_186,FROM_STATE_REG_187,FROM_STATE_REG_188,FROM_STATE_REG_189,FROM_STATE_REG_190,FROM_STATE_REG_191,FROM_STATE_REG_192,FROM_STATE_REG_193,FROM_STATE_REG_194,FROM_STATE_REG_195,FROM_STATE_REG_196,FROM_STATE_REG_197,FROM_STATE_REG_198,FROM_STATE_REG_199,FROM_STATE_REG_200,FROM_STATE_REG_201,FROM_STATE_REG_202,FROM_STATE_REG_203,FROM_STATE_REG_204,FROM_STATE_REG_205,FROM_STATE_REG_206,FROM_STATE_REG_207,FROM_STATE_REG_208,FROM_STATE_REG_209,FROM_STATE_REG_210,FROM_STATE_REG_211,FROM_STATE_REG_212,FROM_STATE_REG_213,FROM_STATE_REG_214,FROM_STATE_REG_215,FROM_STATE_REG_216,FROM_STATE_REG_217,FROM_STATE_REG_218,FROM_STATE_REG_219,FROM_STATE_REG_220,FROM_STATE_REG_221,FROM_STATE_REG_222,FROM_STATE_REG_223,FROM_STATE_REG_224,FROM_STATE_REG_225,FROM_STATE_REG_226,FROM_STATE_REG_227,FROM_STATE_REG_228,FROM_STATE_REG_229,FROM_STATE_REG_230,FROM_STATE_REG_231,FROM_STATE_REG_232,FROM_STATE_REG_233,FROM_STATE_REG_234,FROM_STATE_REG_235,FROM_STATE_REG_236,FROM_STATE_REG_237,FROM_STATE_REG_238,FROM_STATE_REG_239,FROM_STATE_REG_240,FROM_STATE_REG_241,FROM_STATE_REG_242,FROM_STATE_REG_243,FROM_STATE_REG_244,FROM_STATE_REG_245,FROM_STATE_REG_246,FROM_STATE_REG_247,FROM_STATE_REG_248,FROM_STATE_REG_249,FROM_STATE_REG_250,FROM_STATE_REG_251,FROM_STATE_REG_252,FROM_STATE_REG_253,FROM_STATE_REG_254,FROM_STATE_REG_255,FROM_STATE_REG_256,FROM_STATE_REG_257,FROM_STATE_REG_258,FROM_STATE_REG_259,FROM_STATE_REG_260,FROM_STATE_REG_261,FROM_STATE_REG_262,FROM_STATE_REG_263,FROM_STATE_REG_264,FROM_STATE_REG_265,FROM_STATE_REG_266,FROM_STATE_REG_267,FROM_STATE_REG_268,FROM_STATE_REG_269,FROM_STATE_REG_270,FROM_STATE_REG_271,FROM_STATE_REG_272,FROM_STATE_REG_273,FROM_STATE_REG_274,FROM_STATE_REG_275,FROM_STATE_REG_276,FROM_STATE_REG_277,FROM_STATE_REG_278,FROM_STATE_REG_279,FROM_STATE_REG_280,FROM_STATE_REG_281,FROM_STATE_REG_282,FROM_STATE_REG_283,FROM_STATE_REG_284,FROM_STATE_REG_285,FROM_STATE_REG_286,FROM_STATE_REG_287,FROM_STATE_REG_288,FROM_STATE_REG_289,FROM_STATE_REG_290,FROM_STATE_REG_291,FROM_STATE_REG_292,FROM_STATE_REG_293,FROM_STATE_REG_294,FROM_STATE_REG_295,FROM_STATE_REG_296,FROM_STATE_REG_297,FROM_STATE_REG_298,FROM_STATE_REG_299,FROM_STATE_REG_300,FROM_STATE_REG_301,FROM_STATE_REG_302,FROM_STATE_REG_303,FROM_STATE_REG_304,FROM_STATE_REG_305,FROM_STATE_REG_306,FROM_STATE_REG_307,FROM_STATE_REG_308,FROM_STATE_REG_309,FROM_STATE_REG_310,FROM_STATE_REG_311,FROM_STATE_REG_312,FROM_STATE_REG_313,FROM_STATE_REG_314,FROM_STATE_REG_315,FROM_STATE_REG_316,FROM_STATE_REG_317,FROM_STATE_REG_318,FROM_STATE_REG_319,FROM_STATE_REG_320,FROM_STATE_REG_321,FROM_STATE_REG_322,FROM_STATE_REG_323,FROM_STATE_REG_324,FROM_STATE_REG_325,FROM_STATE_REG_326,FROM_STATE_REG_327,FROM_STATE_REG_328,FROM_STATE_REG_329,FROM_STATE_REG_330,FROM_STATE_REG_331,FROM_STATE_REG_332,FROM_STATE_REG_333,FROM_STATE_REG_334,FROM_STATE_REG_335,FROM_STATE_REG_336,FROM_STATE_REG_337,FROM_STATE_REG_338,FROM_STATE_REG_339,FROM_STATE_REG_340,FROM_STATE_REG_341,FROM_STATE_REG_342,FROM_STATE_REG_343,FROM_STATE_REG_344,FROM_STATE_REG_345,FROM_STATE_REG_346,FROM_STATE_REG_347,FROM_STATE_REG_348,FROM_STATE_REG_349,FROM_STATE_REG_350,FROM_STATE_REG_351,FROM_STATE_REG_352,FROM_STATE_REG_353,FROM_STATE_REG_354,FROM_STATE_REG_355,FROM_STATE_REG_356,FROM_STATE_REG_357,FROM_STATE_REG_358,FROM_STATE_REG_359,FROM_STATE_REG_360,FROM_STATE_REG_361,FROM_STATE_REG_362,FROM_STATE_REG_363,FROM_STATE_REG_364,FROM_STATE_REG_365,FROM_STATE_REG_366,FROM_STATE_REG_367,FROM_STATE_REG_368,FROM_STATE_REG_369,FROM_STATE_REG_370,FROM_STATE_REG_371,FROM_STATE_REG_372,FROM_STATE_REG_373,FROM_STATE_REG_374,FROM_STATE_REG_375,FROM_STATE_REG_376,FROM_STATE_REG_377,FROM_STATE_REG_378,FROM_STATE_REG_379,FROM_STATE_REG_380,FROM_STATE_REG_381,FROM_STATE_REG_382,FROM_STATE_REG_383,FROM_STATE_REG_384,FROM_STATE_REG_385,FROM_STATE_REG_386,FROM_STATE_REG_387,FROM_STATE_REG_388,FROM_STATE_REG_389,FROM_STATE_REG_390,FROM_STATE_REG_391,FROM_STATE_REG_392,FROM_STATE_REG_393,FROM_STATE_REG_394,FROM_STATE_REG_395,FROM_STATE_REG_396,FROM_STATE_REG_397,FROM_STATE_REG_398,FROM_STATE_REG_399,FROM_STATE_REG_400,FROM_STATE_REG_401,FROM_STATE_REG_402,FROM_STATE_REG_403,FROM_STATE_REG_404,FROM_STATE_REG_405,FROM_STATE_REG_406,FROM_STATE_REG_407,FROM_STATE_REG_408,FROM_STATE_REG_409,FROM_STATE_REG_410,FROM_STATE_REG_411,FROM_STATE_REG_412,FROM_STATE_REG_413,FROM_STATE_REG_414,FROM_STATE_REG_415,FROM_STATE_REG_416,FROM_STATE_REG_417,FROM_STATE_REG_418,FROM_STATE_REG_419,FROM_STATE_REG_420,FROM_STATE_REG_421,FROM_STATE_REG_422,FROM_STATE_REG_423,FROM_STATE_REG_424,FROM_STATE_REG_425,FROM_STATE_REG_426,FROM_STATE_REG_427,FROM_STATE_REG_428,FROM_STATE_REG_429,FROM_STATE_REG_430,FROM_STATE_REG_431,FROM_STATE_REG_432,FROM_STATE_REG_433,FROM_STATE_REG_434,FROM_STATE_REG_435,FROM_STATE_REG_436,FROM_STATE_REG_437,FROM_STATE_REG_438,FROM_STATE_REG_439,FROM_STATE_REG_440,FROM_STATE_REG_441,FROM_STATE_REG_442,FROM_STATE_REG_443,FROM_STATE_REG_444,FROM_STATE_REG_445,FROM_STATE_REG_446,FROM_STATE_REG_447,FROM_STATE_REG_448,FROM_STATE_REG_449,FROM_STATE_REG_450,FROM_STATE_REG_451,FROM_STATE_REG_452,FROM_STATE_REG_453,FROM_STATE_REG_454,FROM_STATE_REG_455,FROM_STATE_REG_456,FROM_STATE_REG_457,FROM_STATE_REG_458,FROM_STATE_REG_459,FROM_STATE_REG_460,FROM_STATE_REG_461,FROM_STATE_REG_462,FROM_STATE_REG_463,FROM_STATE_REG_464,FROM_STATE_REG_465,FROM_STATE_REG_466,FROM_STATE_REG_467,FROM_STATE_REG_468,FROM_STATE_REG_469,FROM_STATE_REG_470,FROM_STATE_REG_471,FROM_STATE_REG_472,FROM_STATE_REG_473,FROM_STATE_REG_474,FROM_STATE_REG_475,FROM_STATE_REG_476,FROM_STATE_REG_477,FROM_STATE_REG_478,FROM_STATE_REG_479,FROM_STATE_REG_480,FROM_STATE_REG_481,FROM_STATE_REG_482,FROM_STATE_REG_483,FROM_STATE_REG_484,FROM_STATE_REG_485,FROM_STATE_REG_486,FROM_STATE_REG_487,FROM_STATE_REG_488,FROM_STATE_REG_489,FROM_STATE_REG_490,FROM_STATE_REG_491,FROM_STATE_REG_492,FROM_STATE_REG_493,FROM_STATE_REG_494,FROM_STATE_REG_495,FROM_STATE_REG_496,FROM_STATE_REG_497,FROM_STATE_REG_498,FROM_STATE_REG_499,FROM_STATE_REG_500,FROM_STATE_REG_501,FROM_STATE_REG_502,FROM_STATE_REG_503,FROM_STATE_REG_504,FROM_STATE_REG_505,FROM_STATE_REG_506,FROM_STATE_REG_507,FROM_STATE_REG_508,FROM_STATE_REG_509,FROM_STATE_REG_510,FROM_STATE_REG_511,FROM_STATE_REG_512,FROM_STATE_REG_513,FROM_STATE_REG_514,FROM_STATE_REG_515,FROM_STATE_REG_516,FROM_STATE_REG_517,FROM_STATE_REG_518,FROM_STATE_REG_519,FROM_STATE_REG_520,FROM_STATE_REG_521,FROM_STATE_REG_522,FROM_STATE_REG_523,FROM_STATE_REG_524,FROM_STATE_REG_525,FROM_STATE_REG_526,FROM_STATE_REG_527,FROM_STATE_REG_528,FROM_STATE_REG_529,FROM_STATE_REG_530,FROM_STATE_REG_531,FROM_STATE_REG_532,FROM_STATE_REG_533,FROM_STATE_REG_534,FROM_STATE_REG_535,FROM_STATE_REG_536,FROM_STATE_REG_537,FROM_STATE_REG_538,FROM_STATE_REG_539,FROM_STATE_REG_540,FROM_STATE_REG_541,FROM_STATE_REG_542,FROM_STATE_REG_543,FROM_STATE_REG_544,FROM_STATE_REG_545,FROM_STATE_REG_546,FROM_STATE_REG_547,FROM_STATE_REG_548,FROM_STATE_REG_549,FROM_STATE_REG_550,FROM_STATE_REG_551,FROM_STATE_REG_552,FROM_STATE_REG_553,FROM_STATE_REG_554,FROM_STATE_REG_555,FROM_STATE_REG_556,FROM_STATE_REG_557,FROM_STATE_REG_558,FROM_STATE_REG_559,FROM_STATE_REG_560,FROM_STATE_REG_561,FROM_STATE_REG_562,FROM_STATE_REG_563,FROM_STATE_REG_564,FROM_STATE_REG_565,FROM_STATE_REG_566,FROM_STATE_REG_567,FROM_STATE_REG_568,FROM_STATE_REG_569,FROM_STATE_REG_570,FROM_STATE_REG_571,FROM_STATE_REG_572,FROM_STATE_REG_573,FROM_STATE_REG_574,FROM_STATE_REG_575,FROM_STATE_REG_576,FROM_STATE_REG_577,FROM_STATE_REG_578,FROM_STATE_REG_579,FROM_STATE_REG_580,FROM_STATE_REG_581,FROM_STATE_REG_582,FROM_STATE_REG_583,FROM_STATE_REG_584,FROM_STATE_REG_585,FROM_STATE_REG_586,FROM_STATE_REG_587,FROM_STATE_REG_588,FROM_STATE_REG_589,FROM_STATE_REG_590,FROM_STATE_REG_591,FROM_STATE_REG_592,FROM_STATE_REG_593,FROM_STATE_REG_594,FROM_STATE_REG_595,FROM_STATE_REG_596,FROM_STATE_REG_597,FROM_STATE_REG_598,FROM_STATE_REG_599,FROM_STATE_REG_600,FROM_STATE_REG_601,FROM_STATE_REG_602,FROM_STATE_REG_603,FROM_STATE_REG_604,FROM_STATE_REG_605,FROM_STATE_REG_606,FROM_STATE_REG_607,FROM_STATE_REG_608,FROM_STATE_REG_609,FROM_STATE_REG_610,FROM_STATE_REG_611,FROM_STATE_REG_612,FROM_STATE_REG_613,FROM_STATE_REG_614,FROM_STATE_REG_615,FROM_STATE_REG_616,FROM_STATE_REG_617,FROM_STATE_REG_618,FROM_STATE_REG_619,FROM_STATE_REG_620,FROM_STATE_REG_621,FROM_STATE_REG_622,FROM_STATE_REG_623,FROM_STATE_REG_624,FROM_STATE_REG_625,FROM_STATE_REG_626,FROM_STATE_REG_627,FROM_STATE_REG_628,FROM_STATE_REG_629,FROM_STATE_REG_630,FROM_STATE_REG_631,FROM_STATE_REG_632,FROM_STATE_REG_633,FROM_STATE_REG_634,FROM_STATE_REG_635,FROM_STATE_REG_636,FROM_STATE_REG_637,FROM_STATE_REG_638,FROM_STATE_REG_639,FROM_STATE_REG_640,FROM_STATE_REG_641,FROM_STATE_REG_642,FROM_STATE_REG_643,FROM_STATE_REG_644,FROM_STATE_REG_645,FROM_STATE_REG_646,FROM_STATE_REG_647,FROM_STATE_REG_648,FROM_STATE_REG_649,FROM_STATE_REG_650,FROM_STATE_REG_651,FROM_STATE_REG_652,FROM_STATE_REG_653,FROM_STATE_REG_654,FROM_STATE_REG_655,FROM_STATE_REG_656,FROM_STATE_REG_657,FROM_STATE_REG_658,FROM_STATE_REG_659,FROM_STATE_REG_660,FROM_STATE_REG_661,FROM_STATE_REG_662,FROM_STATE_REG_663,FROM_STATE_REG_664,FROM_STATE_REG_665,FROM_STATE_REG_666,FROM_STATE_REG_667,FROM_STATE_REG_668,FROM_STATE_REG_669,FROM_STATE_REG_670,FROM_STATE_REG_671,FROM_STATE_REG_672,FROM_STATE_REG_673,FROM_STATE_REG_674,FROM_STATE_REG_675,FROM_STATE_REG_676,FROM_STATE_REG_677,FROM_STATE_REG_678,FROM_STATE_REG_679,FROM_STATE_REG_680,FROM_STATE_REG_681,FROM_STATE_REG_682,FROM_STATE_REG_683,FROM_STATE_REG_684,FROM_STATE_REG_685,FROM_STATE_REG_686,FROM_STATE_REG_687,FROM_STATE_REG_688,FROM_STATE_REG_689,FROM_STATE_REG_690,FROM_STATE_REG_691,FROM_STATE_REG_692,FROM_STATE_REG_693,FROM_STATE_REG_694,FROM_STATE_REG_695,FROM_STATE_REG_696,FROM_STATE_REG_697,FROM_STATE_REG_698,FROM_STATE_REG_699,FROM_STATE_REG_700,FROM_STATE_REG_701,FROM_STATE_REG_702,FROM_STATE_REG_703,FROM_STATE_REG_704,FROM_STATE_REG_705,FROM_STATE_REG_706,FROM_STATE_REG_707,FROM_STATE_REG_708,FROM_STATE_REG_709,FROM_STATE_REG_710,FROM_STATE_REG_711,FROM_STATE_REG_712,FROM_STATE_REG_713,FROM_STATE_REG_714,FROM_STATE_REG_715,FROM_STATE_REG_716,FROM_STATE_REG_717,FROM_STATE_REG_718,FROM_STATE_REG_719,FROM_STATE_REG_720,FROM_STATE_REG_721,FROM_STATE_REG_722,FROM_STATE_REG_723,FROM_STATE_REG_724,FROM_STATE_REG_725,FROM_STATE_REG_726,FROM_STATE_REG_727,FROM_STATE_REG_728,FROM_STATE_REG_729,FROM_STATE_REG_730,FROM_STATE_REG_731,FROM_STATE_REG_732,FROM_STATE_REG_733,FROM_STATE_REG_734,FROM_STATE_REG_735,FROM_STATE_REG_736,FROM_STATE_REG_737,FROM_STATE_REG_738,FROM_STATE_REG_739,FROM_STATE_REG_740,FROM_STATE_REG_741,FROM_STATE_REG_742,FROM_STATE_REG_743,FROM_STATE_REG_744,FROM_STATE_REG_745,FROM_STATE_REG_746,FROM_STATE_REG_747,FROM_STATE_REG_748,FROM_STATE_REG_749,FROM_STATE_REG_750,FROM_STATE_REG_751,FROM_STATE_REG_752,FROM_STATE_REG_753,FROM_STATE_REG_754,FROM_STATE_REG_755,FROM_STATE_REG_756,FROM_STATE_REG_757,FROM_STATE_REG_758,FROM_STATE_REG_759,FROM_STATE_REG_760,FROM_STATE_REG_761,FROM_STATE_REG_762,FROM_STATE_REG_763,FROM_STATE_REG_764,FROM_STATE_REG_765,FROM_STATE_REG_766,FROM_STATE_REG_767,FROM_STATE_REG_768,FROM_STATE_REG_769,FROM_STATE_REG_770,FROM_STATE_REG_771,FROM_STATE_REG_772,FROM_STATE_REG_773,FROM_STATE_REG_774,FROM_STATE_REG_775,FROM_STATE_REG_776,FROM_STATE_REG_777,FROM_STATE_REG_778,FROM_STATE_REG_779,FROM_STATE_REG_780,FROM_STATE_REG_781,FROM_STATE_REG_782,FROM_STATE_REG_783,FROM_STATE_REG_784,FROM_STATE_REG_785,FROM_STATE_REG_786,FROM_STATE_REG_787,FROM_STATE_REG_788,FROM_STATE_REG_789,FROM_STATE_REG_790,FROM_STATE_REG_791,FROM_STATE_REG_792,FROM_STATE_REG_793,FROM_STATE_REG_794,FROM_STATE_REG_795,FROM_STATE_REG_796,FROM_STATE_REG_797,FROM_STATE_REG_798,FROM_STATE_REG_799,FROM_STATE_REG_800,FROM_STATE_REG_801,FROM_STATE_REG_802,FROM_STATE_REG_803,FROM_STATE_REG_804,FROM_STATE_REG_805,FROM_STATE_REG_806,FROM_STATE_REG_807,FROM_STATE_REG_808,FROM_STATE_REG_809,FROM_STATE_REG_810,FROM_STATE_REG_811,FROM_STATE_REG_812,FROM_STATE_REG_813,FROM_STATE_REG_814,FROM_STATE_REG_815,FROM_STATE_REG_816,FROM_STATE_REG_817,FROM_STATE_REG_818,FROM_STATE_REG_819,FROM_STATE_REG_820,FROM_STATE_REG_821,FROM_STATE_REG_822,FROM_STATE_REG_823,FROM_STATE_REG_824,FROM_STATE_REG_825,FROM_STATE_REG_826,FROM_STATE_REG_827,FROM_STATE_REG_828,FROM_STATE_REG_829,FROM_STATE_REG_830,FROM_STATE_REG_831,FROM_STATE_REG_832,FROM_STATE_REG_833,FROM_STATE_REG_834,FROM_STATE_REG_835,FROM_STATE_REG_836,FROM_STATE_REG_837,FROM_STATE_REG_838,FROM_STATE_REG_839,FROM_STATE_REG_840,FROM_STATE_REG_841,FROM_STATE_REG_842,FROM_STATE_REG_843,FROM_STATE_REG_844,FROM_STATE_REG_845,FROM_STATE_REG_846,FROM_STATE_REG_847,FROM_STATE_REG_848,FROM_STATE_REG_849,FROM_STATE_REG_850,FROM_STATE_REG_851,FROM_STATE_REG_852,FROM_STATE_REG_853,FROM_STATE_REG_854,FROM_STATE_REG_855,FROM_STATE_REG_856,FROM_STATE_REG_857,FROM_STATE_REG_858,FROM_STATE_REG_859,FROM_STATE_REG_860,FROM_STATE_REG_861,FROM_STATE_REG_862,FROM_STATE_REG_863,FROM_STATE_REG_864,FROM_STATE_REG_865,FROM_STATE_REG_866,FROM_STATE_REG_867,FROM_STATE_REG_868,FROM_STATE_REG_869,FROM_STATE_REG_870,FROM_STATE_REG_871,FROM_STATE_REG_872,FROM_STATE_REG_873,FROM_STATE_REG_874,FROM_STATE_REG_875,FROM_STATE_REG_876,FROM_STATE_REG_877,FROM_STATE_REG_878,FROM_STATE_REG_879,FROM_STATE_REG_880,FROM_STATE_REG_881,FROM_STATE_REG_882,FROM_STATE_REG_883,FROM_STATE_REG_884,FROM_STATE_REG_885,FROM_STATE_REG_886,FROM_STATE_REG_887,FROM_STATE_REG_888,FROM_STATE_REG_889,FROM_STATE_REG_890,FROM_STATE_REG_891,FROM_STATE_REG_892,FROM_STATE_REG_893,FROM_STATE_REG_894,FROM_STATE_REG_895,FROM_STATE_REG_896,FROM_STATE_REG_897,FROM_STATE_REG_898,FROM_STATE_REG_899,FROM_STATE_REG_900,FROM_STATE_REG_901,FROM_STATE_REG_902,FROM_STATE_REG_903,FROM_STATE_REG_904,FROM_STATE_REG_905,FROM_STATE_REG_906,FROM_STATE_REG_907,FROM_STATE_REG_908,FROM_STATE_REG_909,FROM_STATE_REG_910,FROM_STATE_REG_911,FROM_STATE_REG_912,FROM_STATE_REG_913,FROM_STATE_REG_914,FROM_STATE_REG_915,FROM_STATE_REG_916,FROM_STATE_REG_917,FROM_STATE_REG_918,FROM_STATE_REG_919,FROM_STATE_REG_920,FROM_STATE_REG_921,FROM_STATE_REG_922,FROM_STATE_REG_923,FROM_STATE_REG_924,FROM_STATE_REG_925,FROM_STATE_REG_926,FROM_STATE_REG_927,FROM_STATE_REG_928,FROM_STATE_REG_929,FROM_STATE_REG_930,FROM_STATE_REG_931,FROM_STATE_REG_932,FROM_STATE_REG_933,FROM_STATE_REG_934,FROM_STATE_REG_935,FROM_STATE_REG_936,FROM_STATE_REG_937,FROM_STATE_REG_938,FROM_STATE_REG_939,FROM_STATE_REG_940,FROM_STATE_REG_941,FROM_STATE_REG_942,FROM_STATE_REG_943,FROM_STATE_REG_944,FROM_STATE_REG_945,FROM_STATE_REG_946,FROM_STATE_REG_947,FROM_STATE_REG_948,FROM_STATE_REG_949,FROM_STATE_REG_950,FROM_STATE_REG_951,FROM_STATE_REG_952,FROM_STATE_REG_953,FROM_STATE_REG_954,FROM_STATE_REG_955,FROM_STATE_REG_956,FROM_STATE_REG_957,FROM_STATE_REG_958,FROM_STATE_REG_959,FROM_STATE_REG_960,FROM_STATE_REG_961,FROM_STATE_REG_962,FROM_STATE_REG_963,FROM_STATE_REG_964,FROM_STATE_REG_965,FROM_STATE_REG_966,FROM_STATE_REG_967,FROM_STATE_REG_968,FROM_STATE_REG_969,FROM_STATE_REG_970,FROM_STATE_REG_971,FROM_STATE_REG_972,FROM_STATE_REG_973,FROM_STATE_REG_974,FROM_STATE_REG_975,FROM_STATE_REG_976,FROM_STATE_REG_977,FROM_STATE_REG_978,FROM_STATE_REG_979,FROM_STATE_REG_980,FROM_STATE_REG_981,FROM_STATE_REG_982,FROM_STATE_REG_983,FROM_STATE_REG_984,FROM_STATE_REG_985,FROM_STATE_REG_986,FROM_STATE_REG_987,FROM_STATE_REG_988,FROM_STATE_REG_989,FROM_STATE_REG_990,FROM_STATE_REG_991,FROM_STATE_REG_992,FROM_STATE_REG_993,FROM_STATE_REG_994,FROM_STATE_REG_995,FROM_STATE_REG_996,FROM_STATE_REG_997,FROM_STATE_REG_998,FROM_STATE_REG_999,FROM_STATE_REG_1000,FROM_STATE_REG_1001,FROM_STATE_REG_1002,FROM_STATE_REG_1003,FROM_STATE_REG_1004,FROM_STATE_REG_1005,FROM_STATE_REG_1006,FROM_STATE_REG_1007,FROM_STATE_REG_1008,FROM_STATE_REG_1009,FROM_STATE_REG_1010,FROM_STATE_REG_1011,FROM_STATE_REG_1012,FROM_STATE_REG_1013,FROM_STATE_REG_1014,FROM_STATE_REG_1015,FROM_STATE_REG_1016,FROM_STATE_REG_1017,FROM_STATE_REG_1018,FROM_STATE_REG_1019,FROM_STATE_REG_1020,FROM_STATE_REG_1021,FROM_STATE_REG_1022,FROM_STATE_REG_1023: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_SELECTION_UNIT_0,FROM_SELECTION_UNIT_1,FROM_SELECTION_UNIT_2,FROM_SELECTION_UNIT_3,FROM_SELECTION_UNIT_4,FROM_SELECTION_UNIT_5,FROM_SELECTION_UNIT_6,FROM_SELECTION_UNIT_7,FROM_SELECTION_UNIT_8,FROM_SELECTION_UNIT_9,FROM_SELECTION_UNIT_10,FROM_SELECTION_UNIT_11,FROM_SELECTION_UNIT_12,FROM_SELECTION_UNIT_13,FROM_SELECTION_UNIT_14,FROM_SELECTION_UNIT_15,FROM_SELECTION_UNIT_16,FROM_SELECTION_UNIT_17,FROM_SELECTION_UNIT_18,FROM_SELECTION_UNIT_19,FROM_SELECTION_UNIT_20,FROM_SELECTION_UNIT_21,FROM_SELECTION_UNIT_22,FROM_SELECTION_UNIT_23,FROM_SELECTION_UNIT_24,FROM_SELECTION_UNIT_25,FROM_SELECTION_UNIT_26,FROM_SELECTION_UNIT_27,FROM_SELECTION_UNIT_28,FROM_SELECTION_UNIT_29,FROM_SELECTION_UNIT_30,FROM_SELECTION_UNIT_31,FROM_SELECTION_UNIT_32,FROM_SELECTION_UNIT_33,FROM_SELECTION_UNIT_34,FROM_SELECTION_UNIT_35,FROM_SELECTION_UNIT_36,FROM_SELECTION_UNIT_37,FROM_SELECTION_UNIT_38,FROM_SELECTION_UNIT_39,FROM_SELECTION_UNIT_40,FROM_SELECTION_UNIT_41,FROM_SELECTION_UNIT_42,FROM_SELECTION_UNIT_43,FROM_SELECTION_UNIT_44,FROM_SELECTION_UNIT_45,FROM_SELECTION_UNIT_46,FROM_SELECTION_UNIT_47,FROM_SELECTION_UNIT_48,FROM_SELECTION_UNIT_49,FROM_SELECTION_UNIT_50,FROM_SELECTION_UNIT_51,FROM_SELECTION_UNIT_52,FROM_SELECTION_UNIT_53,FROM_SELECTION_UNIT_54,FROM_SELECTION_UNIT_55,FROM_SELECTION_UNIT_56,FROM_SELECTION_UNIT_57,FROM_SELECTION_UNIT_58,FROM_SELECTION_UNIT_59,FROM_SELECTION_UNIT_60,FROM_SELECTION_UNIT_61,FROM_SELECTION_UNIT_62,FROM_SELECTION_UNIT_63,FROM_SELECTION_UNIT_64,FROM_SELECTION_UNIT_65,FROM_SELECTION_UNIT_66,FROM_SELECTION_UNIT_67,FROM_SELECTION_UNIT_68,FROM_SELECTION_UNIT_69,FROM_SELECTION_UNIT_70,FROM_SELECTION_UNIT_71,FROM_SELECTION_UNIT_72,FROM_SELECTION_UNIT_73,FROM_SELECTION_UNIT_74,FROM_SELECTION_UNIT_75,FROM_SELECTION_UNIT_76,FROM_SELECTION_UNIT_77,FROM_SELECTION_UNIT_78,FROM_SELECTION_UNIT_79,FROM_SELECTION_UNIT_80,FROM_SELECTION_UNIT_81,FROM_SELECTION_UNIT_82,FROM_SELECTION_UNIT_83,FROM_SELECTION_UNIT_84,FROM_SELECTION_UNIT_85,FROM_SELECTION_UNIT_86,FROM_SELECTION_UNIT_87,FROM_SELECTION_UNIT_88,FROM_SELECTION_UNIT_89,FROM_SELECTION_UNIT_90,FROM_SELECTION_UNIT_91,FROM_SELECTION_UNIT_92,FROM_SELECTION_UNIT_93,FROM_SELECTION_UNIT_94,FROM_SELECTION_UNIT_95,FROM_SELECTION_UNIT_96,FROM_SELECTION_UNIT_97,FROM_SELECTION_UNIT_98,FROM_SELECTION_UNIT_99,FROM_SELECTION_UNIT_100,FROM_SELECTION_UNIT_101,FROM_SELECTION_UNIT_102,FROM_SELECTION_UNIT_103,FROM_SELECTION_UNIT_104,FROM_SELECTION_UNIT_105,FROM_SELECTION_UNIT_106,FROM_SELECTION_UNIT_107,FROM_SELECTION_UNIT_108,FROM_SELECTION_UNIT_109,FROM_SELECTION_UNIT_110,FROM_SELECTION_UNIT_111,FROM_SELECTION_UNIT_112,FROM_SELECTION_UNIT_113,FROM_SELECTION_UNIT_114,FROM_SELECTION_UNIT_115,FROM_SELECTION_UNIT_116,FROM_SELECTION_UNIT_117,FROM_SELECTION_UNIT_118,FROM_SELECTION_UNIT_119,FROM_SELECTION_UNIT_120,FROM_SELECTION_UNIT_121,FROM_SELECTION_UNIT_122,FROM_SELECTION_UNIT_123,FROM_SELECTION_UNIT_124,FROM_SELECTION_UNIT_125,FROM_SELECTION_UNIT_126,FROM_SELECTION_UNIT_127,FROM_SELECTION_UNIT_128,FROM_SELECTION_UNIT_129,FROM_SELECTION_UNIT_130,FROM_SELECTION_UNIT_131,FROM_SELECTION_UNIT_132,FROM_SELECTION_UNIT_133,FROM_SELECTION_UNIT_134,FROM_SELECTION_UNIT_135,FROM_SELECTION_UNIT_136,FROM_SELECTION_UNIT_137,FROM_SELECTION_UNIT_138,FROM_SELECTION_UNIT_139,FROM_SELECTION_UNIT_140,FROM_SELECTION_UNIT_141,FROM_SELECTION_UNIT_142,FROM_SELECTION_UNIT_143,FROM_SELECTION_UNIT_144,FROM_SELECTION_UNIT_145,FROM_SELECTION_UNIT_146,FROM_SELECTION_UNIT_147,FROM_SELECTION_UNIT_148,FROM_SELECTION_UNIT_149,FROM_SELECTION_UNIT_150,FROM_SELECTION_UNIT_151,FROM_SELECTION_UNIT_152,FROM_SELECTION_UNIT_153,FROM_SELECTION_UNIT_154,FROM_SELECTION_UNIT_155,FROM_SELECTION_UNIT_156,FROM_SELECTION_UNIT_157,FROM_SELECTION_UNIT_158,FROM_SELECTION_UNIT_159,FROM_SELECTION_UNIT_160,FROM_SELECTION_UNIT_161,FROM_SELECTION_UNIT_162,FROM_SELECTION_UNIT_163,FROM_SELECTION_UNIT_164,FROM_SELECTION_UNIT_165,FROM_SELECTION_UNIT_166,FROM_SELECTION_UNIT_167,FROM_SELECTION_UNIT_168,FROM_SELECTION_UNIT_169,FROM_SELECTION_UNIT_170,FROM_SELECTION_UNIT_171,FROM_SELECTION_UNIT_172,FROM_SELECTION_UNIT_173,FROM_SELECTION_UNIT_174,FROM_SELECTION_UNIT_175,FROM_SELECTION_UNIT_176,FROM_SELECTION_UNIT_177,FROM_SELECTION_UNIT_178,FROM_SELECTION_UNIT_179,FROM_SELECTION_UNIT_180,FROM_SELECTION_UNIT_181,FROM_SELECTION_UNIT_182,FROM_SELECTION_UNIT_183,FROM_SELECTION_UNIT_184,FROM_SELECTION_UNIT_185,FROM_SELECTION_UNIT_186,FROM_SELECTION_UNIT_187,FROM_SELECTION_UNIT_188,FROM_SELECTION_UNIT_189,FROM_SELECTION_UNIT_190,FROM_SELECTION_UNIT_191,FROM_SELECTION_UNIT_192,FROM_SELECTION_UNIT_193,FROM_SELECTION_UNIT_194,FROM_SELECTION_UNIT_195,FROM_SELECTION_UNIT_196,FROM_SELECTION_UNIT_197,FROM_SELECTION_UNIT_198,FROM_SELECTION_UNIT_199,FROM_SELECTION_UNIT_200,FROM_SELECTION_UNIT_201,FROM_SELECTION_UNIT_202,FROM_SELECTION_UNIT_203,FROM_SELECTION_UNIT_204,FROM_SELECTION_UNIT_205,FROM_SELECTION_UNIT_206,FROM_SELECTION_UNIT_207,FROM_SELECTION_UNIT_208,FROM_SELECTION_UNIT_209,FROM_SELECTION_UNIT_210,FROM_SELECTION_UNIT_211,FROM_SELECTION_UNIT_212,FROM_SELECTION_UNIT_213,FROM_SELECTION_UNIT_214,FROM_SELECTION_UNIT_215,FROM_SELECTION_UNIT_216,FROM_SELECTION_UNIT_217,FROM_SELECTION_UNIT_218,FROM_SELECTION_UNIT_219,FROM_SELECTION_UNIT_220,FROM_SELECTION_UNIT_221,FROM_SELECTION_UNIT_222,FROM_SELECTION_UNIT_223,FROM_SELECTION_UNIT_224,FROM_SELECTION_UNIT_225,FROM_SELECTION_UNIT_226,FROM_SELECTION_UNIT_227,FROM_SELECTION_UNIT_228,FROM_SELECTION_UNIT_229,FROM_SELECTION_UNIT_230,FROM_SELECTION_UNIT_231,FROM_SELECTION_UNIT_232,FROM_SELECTION_UNIT_233,FROM_SELECTION_UNIT_234,FROM_SELECTION_UNIT_235,FROM_SELECTION_UNIT_236,FROM_SELECTION_UNIT_237,FROM_SELECTION_UNIT_238,FROM_SELECTION_UNIT_239,FROM_SELECTION_UNIT_240,FROM_SELECTION_UNIT_241,FROM_SELECTION_UNIT_242,FROM_SELECTION_UNIT_243,FROM_SELECTION_UNIT_244,FROM_SELECTION_UNIT_245,FROM_SELECTION_UNIT_246,FROM_SELECTION_UNIT_247,FROM_SELECTION_UNIT_248,FROM_SELECTION_UNIT_249,FROM_SELECTION_UNIT_250,FROM_SELECTION_UNIT_251,FROM_SELECTION_UNIT_252,FROM_SELECTION_UNIT_253,FROM_SELECTION_UNIT_254,FROM_SELECTION_UNIT_255,FROM_SELECTION_UNIT_256,FROM_SELECTION_UNIT_257,FROM_SELECTION_UNIT_258,FROM_SELECTION_UNIT_259,FROM_SELECTION_UNIT_260,FROM_SELECTION_UNIT_261,FROM_SELECTION_UNIT_262,FROM_SELECTION_UNIT_263,FROM_SELECTION_UNIT_264,FROM_SELECTION_UNIT_265,FROM_SELECTION_UNIT_266,FROM_SELECTION_UNIT_267,FROM_SELECTION_UNIT_268,FROM_SELECTION_UNIT_269,FROM_SELECTION_UNIT_270,FROM_SELECTION_UNIT_271,FROM_SELECTION_UNIT_272,FROM_SELECTION_UNIT_273,FROM_SELECTION_UNIT_274,FROM_SELECTION_UNIT_275,FROM_SELECTION_UNIT_276,FROM_SELECTION_UNIT_277,FROM_SELECTION_UNIT_278,FROM_SELECTION_UNIT_279,FROM_SELECTION_UNIT_280,FROM_SELECTION_UNIT_281,FROM_SELECTION_UNIT_282,FROM_SELECTION_UNIT_283,FROM_SELECTION_UNIT_284,FROM_SELECTION_UNIT_285,FROM_SELECTION_UNIT_286,FROM_SELECTION_UNIT_287,FROM_SELECTION_UNIT_288,FROM_SELECTION_UNIT_289,FROM_SELECTION_UNIT_290,FROM_SELECTION_UNIT_291,FROM_SELECTION_UNIT_292,FROM_SELECTION_UNIT_293,FROM_SELECTION_UNIT_294,FROM_SELECTION_UNIT_295,FROM_SELECTION_UNIT_296,FROM_SELECTION_UNIT_297,FROM_SELECTION_UNIT_298,FROM_SELECTION_UNIT_299,FROM_SELECTION_UNIT_300,FROM_SELECTION_UNIT_301,FROM_SELECTION_UNIT_302,FROM_SELECTION_UNIT_303,FROM_SELECTION_UNIT_304,FROM_SELECTION_UNIT_305,FROM_SELECTION_UNIT_306,FROM_SELECTION_UNIT_307,FROM_SELECTION_UNIT_308,FROM_SELECTION_UNIT_309,FROM_SELECTION_UNIT_310,FROM_SELECTION_UNIT_311,FROM_SELECTION_UNIT_312,FROM_SELECTION_UNIT_313,FROM_SELECTION_UNIT_314,FROM_SELECTION_UNIT_315,FROM_SELECTION_UNIT_316,FROM_SELECTION_UNIT_317,FROM_SELECTION_UNIT_318,FROM_SELECTION_UNIT_319,FROM_SELECTION_UNIT_320,FROM_SELECTION_UNIT_321,FROM_SELECTION_UNIT_322,FROM_SELECTION_UNIT_323,FROM_SELECTION_UNIT_324,FROM_SELECTION_UNIT_325,FROM_SELECTION_UNIT_326,FROM_SELECTION_UNIT_327,FROM_SELECTION_UNIT_328,FROM_SELECTION_UNIT_329,FROM_SELECTION_UNIT_330,FROM_SELECTION_UNIT_331,FROM_SELECTION_UNIT_332,FROM_SELECTION_UNIT_333,FROM_SELECTION_UNIT_334,FROM_SELECTION_UNIT_335,FROM_SELECTION_UNIT_336,FROM_SELECTION_UNIT_337,FROM_SELECTION_UNIT_338,FROM_SELECTION_UNIT_339,FROM_SELECTION_UNIT_340,FROM_SELECTION_UNIT_341,FROM_SELECTION_UNIT_342,FROM_SELECTION_UNIT_343,FROM_SELECTION_UNIT_344,FROM_SELECTION_UNIT_345,FROM_SELECTION_UNIT_346,FROM_SELECTION_UNIT_347,FROM_SELECTION_UNIT_348,FROM_SELECTION_UNIT_349,FROM_SELECTION_UNIT_350,FROM_SELECTION_UNIT_351,FROM_SELECTION_UNIT_352,FROM_SELECTION_UNIT_353,FROM_SELECTION_UNIT_354,FROM_SELECTION_UNIT_355,FROM_SELECTION_UNIT_356,FROM_SELECTION_UNIT_357,FROM_SELECTION_UNIT_358,FROM_SELECTION_UNIT_359,FROM_SELECTION_UNIT_360,FROM_SELECTION_UNIT_361,FROM_SELECTION_UNIT_362,FROM_SELECTION_UNIT_363,FROM_SELECTION_UNIT_364,FROM_SELECTION_UNIT_365,FROM_SELECTION_UNIT_366,FROM_SELECTION_UNIT_367,FROM_SELECTION_UNIT_368,FROM_SELECTION_UNIT_369,FROM_SELECTION_UNIT_370,FROM_SELECTION_UNIT_371,FROM_SELECTION_UNIT_372,FROM_SELECTION_UNIT_373,FROM_SELECTION_UNIT_374,FROM_SELECTION_UNIT_375,FROM_SELECTION_UNIT_376,FROM_SELECTION_UNIT_377,FROM_SELECTION_UNIT_378,FROM_SELECTION_UNIT_379,FROM_SELECTION_UNIT_380,FROM_SELECTION_UNIT_381,FROM_SELECTION_UNIT_382,FROM_SELECTION_UNIT_383,FROM_SELECTION_UNIT_384,FROM_SELECTION_UNIT_385,FROM_SELECTION_UNIT_386,FROM_SELECTION_UNIT_387,FROM_SELECTION_UNIT_388,FROM_SELECTION_UNIT_389,FROM_SELECTION_UNIT_390,FROM_SELECTION_UNIT_391,FROM_SELECTION_UNIT_392,FROM_SELECTION_UNIT_393,FROM_SELECTION_UNIT_394,FROM_SELECTION_UNIT_395,FROM_SELECTION_UNIT_396,FROM_SELECTION_UNIT_397,FROM_SELECTION_UNIT_398,FROM_SELECTION_UNIT_399,FROM_SELECTION_UNIT_400,FROM_SELECTION_UNIT_401,FROM_SELECTION_UNIT_402,FROM_SELECTION_UNIT_403,FROM_SELECTION_UNIT_404,FROM_SELECTION_UNIT_405,FROM_SELECTION_UNIT_406,FROM_SELECTION_UNIT_407,FROM_SELECTION_UNIT_408,FROM_SELECTION_UNIT_409,FROM_SELECTION_UNIT_410,FROM_SELECTION_UNIT_411,FROM_SELECTION_UNIT_412,FROM_SELECTION_UNIT_413,FROM_SELECTION_UNIT_414,FROM_SELECTION_UNIT_415,FROM_SELECTION_UNIT_416,FROM_SELECTION_UNIT_417,FROM_SELECTION_UNIT_418,FROM_SELECTION_UNIT_419,FROM_SELECTION_UNIT_420,FROM_SELECTION_UNIT_421,FROM_SELECTION_UNIT_422,FROM_SELECTION_UNIT_423,FROM_SELECTION_UNIT_424,FROM_SELECTION_UNIT_425,FROM_SELECTION_UNIT_426,FROM_SELECTION_UNIT_427,FROM_SELECTION_UNIT_428,FROM_SELECTION_UNIT_429,FROM_SELECTION_UNIT_430,FROM_SELECTION_UNIT_431,FROM_SELECTION_UNIT_432,FROM_SELECTION_UNIT_433,FROM_SELECTION_UNIT_434,FROM_SELECTION_UNIT_435,FROM_SELECTION_UNIT_436,FROM_SELECTION_UNIT_437,FROM_SELECTION_UNIT_438,FROM_SELECTION_UNIT_439,FROM_SELECTION_UNIT_440,FROM_SELECTION_UNIT_441,FROM_SELECTION_UNIT_442,FROM_SELECTION_UNIT_443,FROM_SELECTION_UNIT_444,FROM_SELECTION_UNIT_445,FROM_SELECTION_UNIT_446,FROM_SELECTION_UNIT_447,FROM_SELECTION_UNIT_448,FROM_SELECTION_UNIT_449,FROM_SELECTION_UNIT_450,FROM_SELECTION_UNIT_451,FROM_SELECTION_UNIT_452,FROM_SELECTION_UNIT_453,FROM_SELECTION_UNIT_454,FROM_SELECTION_UNIT_455,FROM_SELECTION_UNIT_456,FROM_SELECTION_UNIT_457,FROM_SELECTION_UNIT_458,FROM_SELECTION_UNIT_459,FROM_SELECTION_UNIT_460,FROM_SELECTION_UNIT_461,FROM_SELECTION_UNIT_462,FROM_SELECTION_UNIT_463,FROM_SELECTION_UNIT_464,FROM_SELECTION_UNIT_465,FROM_SELECTION_UNIT_466,FROM_SELECTION_UNIT_467,FROM_SELECTION_UNIT_468,FROM_SELECTION_UNIT_469,FROM_SELECTION_UNIT_470,FROM_SELECTION_UNIT_471,FROM_SELECTION_UNIT_472,FROM_SELECTION_UNIT_473,FROM_SELECTION_UNIT_474,FROM_SELECTION_UNIT_475,FROM_SELECTION_UNIT_476,FROM_SELECTION_UNIT_477,FROM_SELECTION_UNIT_478,FROM_SELECTION_UNIT_479,FROM_SELECTION_UNIT_480,FROM_SELECTION_UNIT_481,FROM_SELECTION_UNIT_482,FROM_SELECTION_UNIT_483,FROM_SELECTION_UNIT_484,FROM_SELECTION_UNIT_485,FROM_SELECTION_UNIT_486,FROM_SELECTION_UNIT_487,FROM_SELECTION_UNIT_488,FROM_SELECTION_UNIT_489,FROM_SELECTION_UNIT_490,FROM_SELECTION_UNIT_491,FROM_SELECTION_UNIT_492,FROM_SELECTION_UNIT_493,FROM_SELECTION_UNIT_494,FROM_SELECTION_UNIT_495,FROM_SELECTION_UNIT_496,FROM_SELECTION_UNIT_497,FROM_SELECTION_UNIT_498,FROM_SELECTION_UNIT_499,FROM_SELECTION_UNIT_500,FROM_SELECTION_UNIT_501,FROM_SELECTION_UNIT_502,FROM_SELECTION_UNIT_503,FROM_SELECTION_UNIT_504,FROM_SELECTION_UNIT_505,FROM_SELECTION_UNIT_506,FROM_SELECTION_UNIT_507,FROM_SELECTION_UNIT_508,FROM_SELECTION_UNIT_509,FROM_SELECTION_UNIT_510,FROM_SELECTION_UNIT_511,FROM_SELECTION_UNIT_512,FROM_SELECTION_UNIT_513,FROM_SELECTION_UNIT_514,FROM_SELECTION_UNIT_515,FROM_SELECTION_UNIT_516,FROM_SELECTION_UNIT_517,FROM_SELECTION_UNIT_518,FROM_SELECTION_UNIT_519,FROM_SELECTION_UNIT_520,FROM_SELECTION_UNIT_521,FROM_SELECTION_UNIT_522,FROM_SELECTION_UNIT_523,FROM_SELECTION_UNIT_524,FROM_SELECTION_UNIT_525,FROM_SELECTION_UNIT_526,FROM_SELECTION_UNIT_527,FROM_SELECTION_UNIT_528,FROM_SELECTION_UNIT_529,FROM_SELECTION_UNIT_530,FROM_SELECTION_UNIT_531,FROM_SELECTION_UNIT_532,FROM_SELECTION_UNIT_533,FROM_SELECTION_UNIT_534,FROM_SELECTION_UNIT_535,FROM_SELECTION_UNIT_536,FROM_SELECTION_UNIT_537,FROM_SELECTION_UNIT_538,FROM_SELECTION_UNIT_539,FROM_SELECTION_UNIT_540,FROM_SELECTION_UNIT_541,FROM_SELECTION_UNIT_542,FROM_SELECTION_UNIT_543,FROM_SELECTION_UNIT_544,FROM_SELECTION_UNIT_545,FROM_SELECTION_UNIT_546,FROM_SELECTION_UNIT_547,FROM_SELECTION_UNIT_548,FROM_SELECTION_UNIT_549,FROM_SELECTION_UNIT_550,FROM_SELECTION_UNIT_551,FROM_SELECTION_UNIT_552,FROM_SELECTION_UNIT_553,FROM_SELECTION_UNIT_554,FROM_SELECTION_UNIT_555,FROM_SELECTION_UNIT_556,FROM_SELECTION_UNIT_557,FROM_SELECTION_UNIT_558,FROM_SELECTION_UNIT_559,FROM_SELECTION_UNIT_560,FROM_SELECTION_UNIT_561,FROM_SELECTION_UNIT_562,FROM_SELECTION_UNIT_563,FROM_SELECTION_UNIT_564,FROM_SELECTION_UNIT_565,FROM_SELECTION_UNIT_566,FROM_SELECTION_UNIT_567,FROM_SELECTION_UNIT_568,FROM_SELECTION_UNIT_569,FROM_SELECTION_UNIT_570,FROM_SELECTION_UNIT_571,FROM_SELECTION_UNIT_572,FROM_SELECTION_UNIT_573,FROM_SELECTION_UNIT_574,FROM_SELECTION_UNIT_575,FROM_SELECTION_UNIT_576,FROM_SELECTION_UNIT_577,FROM_SELECTION_UNIT_578,FROM_SELECTION_UNIT_579,FROM_SELECTION_UNIT_580,FROM_SELECTION_UNIT_581,FROM_SELECTION_UNIT_582,FROM_SELECTION_UNIT_583,FROM_SELECTION_UNIT_584,FROM_SELECTION_UNIT_585,FROM_SELECTION_UNIT_586,FROM_SELECTION_UNIT_587,FROM_SELECTION_UNIT_588,FROM_SELECTION_UNIT_589,FROM_SELECTION_UNIT_590,FROM_SELECTION_UNIT_591,FROM_SELECTION_UNIT_592,FROM_SELECTION_UNIT_593,FROM_SELECTION_UNIT_594,FROM_SELECTION_UNIT_595,FROM_SELECTION_UNIT_596,FROM_SELECTION_UNIT_597,FROM_SELECTION_UNIT_598,FROM_SELECTION_UNIT_599,FROM_SELECTION_UNIT_600,FROM_SELECTION_UNIT_601,FROM_SELECTION_UNIT_602,FROM_SELECTION_UNIT_603,FROM_SELECTION_UNIT_604,FROM_SELECTION_UNIT_605,FROM_SELECTION_UNIT_606,FROM_SELECTION_UNIT_607,FROM_SELECTION_UNIT_608,FROM_SELECTION_UNIT_609,FROM_SELECTION_UNIT_610,FROM_SELECTION_UNIT_611,FROM_SELECTION_UNIT_612,FROM_SELECTION_UNIT_613,FROM_SELECTION_UNIT_614,FROM_SELECTION_UNIT_615,FROM_SELECTION_UNIT_616,FROM_SELECTION_UNIT_617,FROM_SELECTION_UNIT_618,FROM_SELECTION_UNIT_619,FROM_SELECTION_UNIT_620,FROM_SELECTION_UNIT_621,FROM_SELECTION_UNIT_622,FROM_SELECTION_UNIT_623,FROM_SELECTION_UNIT_624,FROM_SELECTION_UNIT_625,FROM_SELECTION_UNIT_626,FROM_SELECTION_UNIT_627,FROM_SELECTION_UNIT_628,FROM_SELECTION_UNIT_629,FROM_SELECTION_UNIT_630,FROM_SELECTION_UNIT_631,FROM_SELECTION_UNIT_632,FROM_SELECTION_UNIT_633,FROM_SELECTION_UNIT_634,FROM_SELECTION_UNIT_635,FROM_SELECTION_UNIT_636,FROM_SELECTION_UNIT_637,FROM_SELECTION_UNIT_638,FROM_SELECTION_UNIT_639,FROM_SELECTION_UNIT_640,FROM_SELECTION_UNIT_641,FROM_SELECTION_UNIT_642,FROM_SELECTION_UNIT_643,FROM_SELECTION_UNIT_644,FROM_SELECTION_UNIT_645,FROM_SELECTION_UNIT_646,FROM_SELECTION_UNIT_647,FROM_SELECTION_UNIT_648,FROM_SELECTION_UNIT_649,FROM_SELECTION_UNIT_650,FROM_SELECTION_UNIT_651,FROM_SELECTION_UNIT_652,FROM_SELECTION_UNIT_653,FROM_SELECTION_UNIT_654,FROM_SELECTION_UNIT_655,FROM_SELECTION_UNIT_656,FROM_SELECTION_UNIT_657,FROM_SELECTION_UNIT_658,FROM_SELECTION_UNIT_659,FROM_SELECTION_UNIT_660,FROM_SELECTION_UNIT_661,FROM_SELECTION_UNIT_662,FROM_SELECTION_UNIT_663,FROM_SELECTION_UNIT_664,FROM_SELECTION_UNIT_665,FROM_SELECTION_UNIT_666,FROM_SELECTION_UNIT_667,FROM_SELECTION_UNIT_668,FROM_SELECTION_UNIT_669,FROM_SELECTION_UNIT_670,FROM_SELECTION_UNIT_671,FROM_SELECTION_UNIT_672,FROM_SELECTION_UNIT_673,FROM_SELECTION_UNIT_674,FROM_SELECTION_UNIT_675,FROM_SELECTION_UNIT_676,FROM_SELECTION_UNIT_677,FROM_SELECTION_UNIT_678,FROM_SELECTION_UNIT_679,FROM_SELECTION_UNIT_680,FROM_SELECTION_UNIT_681,FROM_SELECTION_UNIT_682,FROM_SELECTION_UNIT_683,FROM_SELECTION_UNIT_684,FROM_SELECTION_UNIT_685,FROM_SELECTION_UNIT_686,FROM_SELECTION_UNIT_687,FROM_SELECTION_UNIT_688,FROM_SELECTION_UNIT_689,FROM_SELECTION_UNIT_690,FROM_SELECTION_UNIT_691,FROM_SELECTION_UNIT_692,FROM_SELECTION_UNIT_693,FROM_SELECTION_UNIT_694,FROM_SELECTION_UNIT_695,FROM_SELECTION_UNIT_696,FROM_SELECTION_UNIT_697,FROM_SELECTION_UNIT_698,FROM_SELECTION_UNIT_699,FROM_SELECTION_UNIT_700,FROM_SELECTION_UNIT_701,FROM_SELECTION_UNIT_702,FROM_SELECTION_UNIT_703,FROM_SELECTION_UNIT_704,FROM_SELECTION_UNIT_705,FROM_SELECTION_UNIT_706,FROM_SELECTION_UNIT_707,FROM_SELECTION_UNIT_708,FROM_SELECTION_UNIT_709,FROM_SELECTION_UNIT_710,FROM_SELECTION_UNIT_711,FROM_SELECTION_UNIT_712,FROM_SELECTION_UNIT_713,FROM_SELECTION_UNIT_714,FROM_SELECTION_UNIT_715,FROM_SELECTION_UNIT_716,FROM_SELECTION_UNIT_717,FROM_SELECTION_UNIT_718,FROM_SELECTION_UNIT_719,FROM_SELECTION_UNIT_720,FROM_SELECTION_UNIT_721,FROM_SELECTION_UNIT_722,FROM_SELECTION_UNIT_723,FROM_SELECTION_UNIT_724,FROM_SELECTION_UNIT_725,FROM_SELECTION_UNIT_726,FROM_SELECTION_UNIT_727,FROM_SELECTION_UNIT_728,FROM_SELECTION_UNIT_729,FROM_SELECTION_UNIT_730,FROM_SELECTION_UNIT_731,FROM_SELECTION_UNIT_732,FROM_SELECTION_UNIT_733,FROM_SELECTION_UNIT_734,FROM_SELECTION_UNIT_735,FROM_SELECTION_UNIT_736,FROM_SELECTION_UNIT_737,FROM_SELECTION_UNIT_738,FROM_SELECTION_UNIT_739,FROM_SELECTION_UNIT_740,FROM_SELECTION_UNIT_741,FROM_SELECTION_UNIT_742,FROM_SELECTION_UNIT_743,FROM_SELECTION_UNIT_744,FROM_SELECTION_UNIT_745,FROM_SELECTION_UNIT_746,FROM_SELECTION_UNIT_747,FROM_SELECTION_UNIT_748,FROM_SELECTION_UNIT_749,FROM_SELECTION_UNIT_750,FROM_SELECTION_UNIT_751,FROM_SELECTION_UNIT_752,FROM_SELECTION_UNIT_753,FROM_SELECTION_UNIT_754,FROM_SELECTION_UNIT_755,FROM_SELECTION_UNIT_756,FROM_SELECTION_UNIT_757,FROM_SELECTION_UNIT_758,FROM_SELECTION_UNIT_759,FROM_SELECTION_UNIT_760,FROM_SELECTION_UNIT_761,FROM_SELECTION_UNIT_762,FROM_SELECTION_UNIT_763,FROM_SELECTION_UNIT_764,FROM_SELECTION_UNIT_765,FROM_SELECTION_UNIT_766,FROM_SELECTION_UNIT_767,FROM_SELECTION_UNIT_768,FROM_SELECTION_UNIT_769,FROM_SELECTION_UNIT_770,FROM_SELECTION_UNIT_771,FROM_SELECTION_UNIT_772,FROM_SELECTION_UNIT_773,FROM_SELECTION_UNIT_774,FROM_SELECTION_UNIT_775,FROM_SELECTION_UNIT_776,FROM_SELECTION_UNIT_777,FROM_SELECTION_UNIT_778,FROM_SELECTION_UNIT_779,FROM_SELECTION_UNIT_780,FROM_SELECTION_UNIT_781,FROM_SELECTION_UNIT_782,FROM_SELECTION_UNIT_783,FROM_SELECTION_UNIT_784,FROM_SELECTION_UNIT_785,FROM_SELECTION_UNIT_786,FROM_SELECTION_UNIT_787,FROM_SELECTION_UNIT_788,FROM_SELECTION_UNIT_789,FROM_SELECTION_UNIT_790,FROM_SELECTION_UNIT_791,FROM_SELECTION_UNIT_792,FROM_SELECTION_UNIT_793,FROM_SELECTION_UNIT_794,FROM_SELECTION_UNIT_795,FROM_SELECTION_UNIT_796,FROM_SELECTION_UNIT_797,FROM_SELECTION_UNIT_798,FROM_SELECTION_UNIT_799,FROM_SELECTION_UNIT_800,FROM_SELECTION_UNIT_801,FROM_SELECTION_UNIT_802,FROM_SELECTION_UNIT_803,FROM_SELECTION_UNIT_804,FROM_SELECTION_UNIT_805,FROM_SELECTION_UNIT_806,FROM_SELECTION_UNIT_807,FROM_SELECTION_UNIT_808,FROM_SELECTION_UNIT_809,FROM_SELECTION_UNIT_810,FROM_SELECTION_UNIT_811,FROM_SELECTION_UNIT_812,FROM_SELECTION_UNIT_813,FROM_SELECTION_UNIT_814,FROM_SELECTION_UNIT_815,FROM_SELECTION_UNIT_816,FROM_SELECTION_UNIT_817,FROM_SELECTION_UNIT_818,FROM_SELECTION_UNIT_819,FROM_SELECTION_UNIT_820,FROM_SELECTION_UNIT_821,FROM_SELECTION_UNIT_822,FROM_SELECTION_UNIT_823,FROM_SELECTION_UNIT_824,FROM_SELECTION_UNIT_825,FROM_SELECTION_UNIT_826,FROM_SELECTION_UNIT_827,FROM_SELECTION_UNIT_828,FROM_SELECTION_UNIT_829,FROM_SELECTION_UNIT_830,FROM_SELECTION_UNIT_831,FROM_SELECTION_UNIT_832,FROM_SELECTION_UNIT_833,FROM_SELECTION_UNIT_834,FROM_SELECTION_UNIT_835,FROM_SELECTION_UNIT_836,FROM_SELECTION_UNIT_837,FROM_SELECTION_UNIT_838,FROM_SELECTION_UNIT_839,FROM_SELECTION_UNIT_840,FROM_SELECTION_UNIT_841,FROM_SELECTION_UNIT_842,FROM_SELECTION_UNIT_843,FROM_SELECTION_UNIT_844,FROM_SELECTION_UNIT_845,FROM_SELECTION_UNIT_846,FROM_SELECTION_UNIT_847,FROM_SELECTION_UNIT_848,FROM_SELECTION_UNIT_849,FROM_SELECTION_UNIT_850,FROM_SELECTION_UNIT_851,FROM_SELECTION_UNIT_852,FROM_SELECTION_UNIT_853,FROM_SELECTION_UNIT_854,FROM_SELECTION_UNIT_855,FROM_SELECTION_UNIT_856,FROM_SELECTION_UNIT_857,FROM_SELECTION_UNIT_858,FROM_SELECTION_UNIT_859,FROM_SELECTION_UNIT_860,FROM_SELECTION_UNIT_861,FROM_SELECTION_UNIT_862,FROM_SELECTION_UNIT_863,FROM_SELECTION_UNIT_864,FROM_SELECTION_UNIT_865,FROM_SELECTION_UNIT_866,FROM_SELECTION_UNIT_867,FROM_SELECTION_UNIT_868,FROM_SELECTION_UNIT_869,FROM_SELECTION_UNIT_870,FROM_SELECTION_UNIT_871,FROM_SELECTION_UNIT_872,FROM_SELECTION_UNIT_873,FROM_SELECTION_UNIT_874,FROM_SELECTION_UNIT_875,FROM_SELECTION_UNIT_876,FROM_SELECTION_UNIT_877,FROM_SELECTION_UNIT_878,FROM_SELECTION_UNIT_879,FROM_SELECTION_UNIT_880,FROM_SELECTION_UNIT_881,FROM_SELECTION_UNIT_882,FROM_SELECTION_UNIT_883,FROM_SELECTION_UNIT_884,FROM_SELECTION_UNIT_885,FROM_SELECTION_UNIT_886,FROM_SELECTION_UNIT_887,FROM_SELECTION_UNIT_888,FROM_SELECTION_UNIT_889,FROM_SELECTION_UNIT_890,FROM_SELECTION_UNIT_891,FROM_SELECTION_UNIT_892,FROM_SELECTION_UNIT_893,FROM_SELECTION_UNIT_894,FROM_SELECTION_UNIT_895,FROM_SELECTION_UNIT_896,FROM_SELECTION_UNIT_897,FROM_SELECTION_UNIT_898,FROM_SELECTION_UNIT_899,FROM_SELECTION_UNIT_900,FROM_SELECTION_UNIT_901,FROM_SELECTION_UNIT_902,FROM_SELECTION_UNIT_903,FROM_SELECTION_UNIT_904,FROM_SELECTION_UNIT_905,FROM_SELECTION_UNIT_906,FROM_SELECTION_UNIT_907,FROM_SELECTION_UNIT_908,FROM_SELECTION_UNIT_909,FROM_SELECTION_UNIT_910,FROM_SELECTION_UNIT_911,FROM_SELECTION_UNIT_912,FROM_SELECTION_UNIT_913,FROM_SELECTION_UNIT_914,FROM_SELECTION_UNIT_915,FROM_SELECTION_UNIT_916,FROM_SELECTION_UNIT_917,FROM_SELECTION_UNIT_918,FROM_SELECTION_UNIT_919,FROM_SELECTION_UNIT_920,FROM_SELECTION_UNIT_921,FROM_SELECTION_UNIT_922,FROM_SELECTION_UNIT_923,FROM_SELECTION_UNIT_924,FROM_SELECTION_UNIT_925,FROM_SELECTION_UNIT_926,FROM_SELECTION_UNIT_927,FROM_SELECTION_UNIT_928,FROM_SELECTION_UNIT_929,FROM_SELECTION_UNIT_930,FROM_SELECTION_UNIT_931,FROM_SELECTION_UNIT_932,FROM_SELECTION_UNIT_933,FROM_SELECTION_UNIT_934,FROM_SELECTION_UNIT_935,FROM_SELECTION_UNIT_936,FROM_SELECTION_UNIT_937,FROM_SELECTION_UNIT_938,FROM_SELECTION_UNIT_939,FROM_SELECTION_UNIT_940,FROM_SELECTION_UNIT_941,FROM_SELECTION_UNIT_942,FROM_SELECTION_UNIT_943,FROM_SELECTION_UNIT_944,FROM_SELECTION_UNIT_945,FROM_SELECTION_UNIT_946,FROM_SELECTION_UNIT_947,FROM_SELECTION_UNIT_948,FROM_SELECTION_UNIT_949,FROM_SELECTION_UNIT_950,FROM_SELECTION_UNIT_951,FROM_SELECTION_UNIT_952,FROM_SELECTION_UNIT_953,FROM_SELECTION_UNIT_954,FROM_SELECTION_UNIT_955,FROM_SELECTION_UNIT_956,FROM_SELECTION_UNIT_957,FROM_SELECTION_UNIT_958,FROM_SELECTION_UNIT_959,FROM_SELECTION_UNIT_960,FROM_SELECTION_UNIT_961,FROM_SELECTION_UNIT_962,FROM_SELECTION_UNIT_963,FROM_SELECTION_UNIT_964,FROM_SELECTION_UNIT_965,FROM_SELECTION_UNIT_966,FROM_SELECTION_UNIT_967,FROM_SELECTION_UNIT_968,FROM_SELECTION_UNIT_969,FROM_SELECTION_UNIT_970,FROM_SELECTION_UNIT_971,FROM_SELECTION_UNIT_972,FROM_SELECTION_UNIT_973,FROM_SELECTION_UNIT_974,FROM_SELECTION_UNIT_975,FROM_SELECTION_UNIT_976,FROM_SELECTION_UNIT_977,FROM_SELECTION_UNIT_978,FROM_SELECTION_UNIT_979,FROM_SELECTION_UNIT_980,FROM_SELECTION_UNIT_981,FROM_SELECTION_UNIT_982,FROM_SELECTION_UNIT_983,FROM_SELECTION_UNIT_984,FROM_SELECTION_UNIT_985,FROM_SELECTION_UNIT_986,FROM_SELECTION_UNIT_987,FROM_SELECTION_UNIT_988,FROM_SELECTION_UNIT_989,FROM_SELECTION_UNIT_990,FROM_SELECTION_UNIT_991,FROM_SELECTION_UNIT_992,FROM_SELECTION_UNIT_993,FROM_SELECTION_UNIT_994,FROM_SELECTION_UNIT_995,FROM_SELECTION_UNIT_996,FROM_SELECTION_UNIT_997,FROM_SELECTION_UNIT_998,FROM_SELECTION_UNIT_999,FROM_SELECTION_UNIT_1000,FROM_SELECTION_UNIT_1001,FROM_SELECTION_UNIT_1002,FROM_SELECTION_UNIT_1003,FROM_SELECTION_UNIT_1004,FROM_SELECTION_UNIT_1005,FROM_SELECTION_UNIT_1006,FROM_SELECTION_UNIT_1007,FROM_SELECTION_UNIT_1008,FROM_SELECTION_UNIT_1009,FROM_SELECTION_UNIT_1010,FROM_SELECTION_UNIT_1011,FROM_SELECTION_UNIT_1012,FROM_SELECTION_UNIT_1013,FROM_SELECTION_UNIT_1014,FROM_SELECTION_UNIT_1015,FROM_SELECTION_UNIT_1016,FROM_SELECTION_UNIT_1017,FROM_SELECTION_UNIT_1018,FROM_SELECTION_UNIT_1019,FROM_SELECTION_UNIT_1020,FROM_SELECTION_UNIT_1021,FROM_SELECTION_UNIT_1022,FROM_SELECTION_UNIT_1023: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_0,FROM_WINDOW_1,FROM_WINDOW_2,FROM_WINDOW_3,FROM_WINDOW_4,FROM_WINDOW_5,FROM_WINDOW_6,FROM_WINDOW_7,FROM_WINDOW_8,FROM_WINDOW_9,FROM_WINDOW_10,FROM_WINDOW_11,FROM_WINDOW_12,FROM_WINDOW_13,FROM_WINDOW_14,FROM_WINDOW_15,FROM_WINDOW_16,FROM_WINDOW_17,FROM_WINDOW_18,FROM_WINDOW_19,FROM_WINDOW_20,FROM_WINDOW_21,FROM_WINDOW_22,FROM_WINDOW_23,FROM_WINDOW_24,FROM_WINDOW_25,FROM_WINDOW_26,FROM_WINDOW_27,FROM_WINDOW_28,FROM_WINDOW_29,FROM_WINDOW_30,FROM_WINDOW_31,FROM_WINDOW_32,FROM_WINDOW_33,FROM_WINDOW_34,FROM_WINDOW_35,FROM_WINDOW_36,FROM_WINDOW_37,FROM_WINDOW_38,FROM_WINDOW_39,FROM_WINDOW_40,FROM_WINDOW_41,FROM_WINDOW_42,FROM_WINDOW_43,FROM_WINDOW_44,FROM_WINDOW_45,FROM_WINDOW_46,FROM_WINDOW_47,FROM_WINDOW_48,FROM_WINDOW_49,FROM_WINDOW_50,FROM_WINDOW_51,FROM_WINDOW_52,FROM_WINDOW_53,FROM_WINDOW_54,FROM_WINDOW_55,FROM_WINDOW_56,FROM_WINDOW_57,FROM_WINDOW_58,FROM_WINDOW_59,FROM_WINDOW_60,FROM_WINDOW_61,FROM_WINDOW_62,FROM_WINDOW_63,FROM_WINDOW_64,FROM_WINDOW_65,FROM_WINDOW_66,FROM_WINDOW_67,FROM_WINDOW_68,FROM_WINDOW_69,FROM_WINDOW_70,FROM_WINDOW_71,FROM_WINDOW_72,FROM_WINDOW_73,FROM_WINDOW_74,FROM_WINDOW_75,FROM_WINDOW_76,FROM_WINDOW_77,FROM_WINDOW_78,FROM_WINDOW_79,FROM_WINDOW_80,FROM_WINDOW_81,FROM_WINDOW_82,FROM_WINDOW_83,FROM_WINDOW_84,FROM_WINDOW_85,FROM_WINDOW_86,FROM_WINDOW_87,FROM_WINDOW_88,FROM_WINDOW_89,FROM_WINDOW_90,FROM_WINDOW_91,FROM_WINDOW_92,FROM_WINDOW_93,FROM_WINDOW_94,FROM_WINDOW_95,FROM_WINDOW_96,FROM_WINDOW_97,FROM_WINDOW_98,FROM_WINDOW_99,FROM_WINDOW_100,FROM_WINDOW_101,FROM_WINDOW_102,FROM_WINDOW_103,FROM_WINDOW_104,FROM_WINDOW_105,FROM_WINDOW_106,FROM_WINDOW_107,FROM_WINDOW_108,FROM_WINDOW_109,FROM_WINDOW_110,FROM_WINDOW_111,FROM_WINDOW_112,FROM_WINDOW_113,FROM_WINDOW_114,FROM_WINDOW_115,FROM_WINDOW_116,FROM_WINDOW_117,FROM_WINDOW_118,FROM_WINDOW_119,FROM_WINDOW_120,FROM_WINDOW_121,FROM_WINDOW_122,FROM_WINDOW_123,FROM_WINDOW_124,FROM_WINDOW_125,FROM_WINDOW_126,FROM_WINDOW_127,FROM_WINDOW_128,FROM_WINDOW_129,FROM_WINDOW_130,FROM_WINDOW_131,FROM_WINDOW_132,FROM_WINDOW_133,FROM_WINDOW_134,FROM_WINDOW_135,FROM_WINDOW_136,FROM_WINDOW_137,FROM_WINDOW_138,FROM_WINDOW_139,FROM_WINDOW_140,FROM_WINDOW_141,FROM_WINDOW_142,FROM_WINDOW_143,FROM_WINDOW_144,FROM_WINDOW_145,FROM_WINDOW_146,FROM_WINDOW_147,FROM_WINDOW_148,FROM_WINDOW_149,FROM_WINDOW_150,FROM_WINDOW_151,FROM_WINDOW_152,FROM_WINDOW_153,FROM_WINDOW_154,FROM_WINDOW_155,FROM_WINDOW_156,FROM_WINDOW_157,FROM_WINDOW_158,FROM_WINDOW_159,FROM_WINDOW_160,FROM_WINDOW_161,FROM_WINDOW_162,FROM_WINDOW_163,FROM_WINDOW_164,FROM_WINDOW_165,FROM_WINDOW_166,FROM_WINDOW_167,FROM_WINDOW_168,FROM_WINDOW_169,FROM_WINDOW_170,FROM_WINDOW_171,FROM_WINDOW_172,FROM_WINDOW_173,FROM_WINDOW_174,FROM_WINDOW_175,FROM_WINDOW_176,FROM_WINDOW_177,FROM_WINDOW_178,FROM_WINDOW_179,FROM_WINDOW_180,FROM_WINDOW_181,FROM_WINDOW_182,FROM_WINDOW_183,FROM_WINDOW_184,FROM_WINDOW_185,FROM_WINDOW_186,FROM_WINDOW_187,FROM_WINDOW_188,FROM_WINDOW_189,FROM_WINDOW_190,FROM_WINDOW_191,FROM_WINDOW_192,FROM_WINDOW_193,FROM_WINDOW_194,FROM_WINDOW_195,FROM_WINDOW_196,FROM_WINDOW_197,FROM_WINDOW_198,FROM_WINDOW_199,FROM_WINDOW_200,FROM_WINDOW_201,FROM_WINDOW_202,FROM_WINDOW_203,FROM_WINDOW_204,FROM_WINDOW_205,FROM_WINDOW_206,FROM_WINDOW_207,FROM_WINDOW_208,FROM_WINDOW_209,FROM_WINDOW_210,FROM_WINDOW_211,FROM_WINDOW_212,FROM_WINDOW_213,FROM_WINDOW_214,FROM_WINDOW_215,FROM_WINDOW_216,FROM_WINDOW_217,FROM_WINDOW_218,FROM_WINDOW_219,FROM_WINDOW_220,FROM_WINDOW_221,FROM_WINDOW_222,FROM_WINDOW_223,FROM_WINDOW_224,FROM_WINDOW_225,FROM_WINDOW_226,FROM_WINDOW_227,FROM_WINDOW_228,FROM_WINDOW_229,FROM_WINDOW_230,FROM_WINDOW_231,FROM_WINDOW_232,FROM_WINDOW_233,FROM_WINDOW_234,FROM_WINDOW_235,FROM_WINDOW_236,FROM_WINDOW_237,FROM_WINDOW_238,FROM_WINDOW_239,FROM_WINDOW_240,FROM_WINDOW_241,FROM_WINDOW_242,FROM_WINDOW_243,FROM_WINDOW_244,FROM_WINDOW_245,FROM_WINDOW_246,FROM_WINDOW_247,FROM_WINDOW_248,FROM_WINDOW_249,FROM_WINDOW_250,FROM_WINDOW_251,FROM_WINDOW_252,FROM_WINDOW_253,FROM_WINDOW_254,FROM_WINDOW_255,FROM_WINDOW_256,FROM_WINDOW_257,FROM_WINDOW_258,FROM_WINDOW_259,FROM_WINDOW_260,FROM_WINDOW_261,FROM_WINDOW_262,FROM_WINDOW_263,FROM_WINDOW_264,FROM_WINDOW_265,FROM_WINDOW_266,FROM_WINDOW_267,FROM_WINDOW_268,FROM_WINDOW_269,FROM_WINDOW_270,FROM_WINDOW_271,FROM_WINDOW_272,FROM_WINDOW_273,FROM_WINDOW_274,FROM_WINDOW_275,FROM_WINDOW_276,FROM_WINDOW_277,FROM_WINDOW_278,FROM_WINDOW_279,FROM_WINDOW_280,FROM_WINDOW_281,FROM_WINDOW_282,FROM_WINDOW_283,FROM_WINDOW_284,FROM_WINDOW_285,FROM_WINDOW_286,FROM_WINDOW_287,FROM_WINDOW_288,FROM_WINDOW_289,FROM_WINDOW_290,FROM_WINDOW_291,FROM_WINDOW_292,FROM_WINDOW_293,FROM_WINDOW_294,FROM_WINDOW_295,FROM_WINDOW_296,FROM_WINDOW_297,FROM_WINDOW_298,FROM_WINDOW_299,FROM_WINDOW_300,FROM_WINDOW_301,FROM_WINDOW_302,FROM_WINDOW_303,FROM_WINDOW_304,FROM_WINDOW_305,FROM_WINDOW_306,FROM_WINDOW_307,FROM_WINDOW_308,FROM_WINDOW_309,FROM_WINDOW_310,FROM_WINDOW_311,FROM_WINDOW_312,FROM_WINDOW_313,FROM_WINDOW_314,FROM_WINDOW_315,FROM_WINDOW_316,FROM_WINDOW_317,FROM_WINDOW_318,FROM_WINDOW_319,FROM_WINDOW_320,FROM_WINDOW_321,FROM_WINDOW_322,FROM_WINDOW_323,FROM_WINDOW_324,FROM_WINDOW_325,FROM_WINDOW_326,FROM_WINDOW_327,FROM_WINDOW_328,FROM_WINDOW_329,FROM_WINDOW_330,FROM_WINDOW_331,FROM_WINDOW_332,FROM_WINDOW_333,FROM_WINDOW_334,FROM_WINDOW_335,FROM_WINDOW_336,FROM_WINDOW_337,FROM_WINDOW_338,FROM_WINDOW_339,FROM_WINDOW_340,FROM_WINDOW_341,FROM_WINDOW_342,FROM_WINDOW_343,FROM_WINDOW_344,FROM_WINDOW_345,FROM_WINDOW_346,FROM_WINDOW_347,FROM_WINDOW_348,FROM_WINDOW_349,FROM_WINDOW_350,FROM_WINDOW_351,FROM_WINDOW_352,FROM_WINDOW_353,FROM_WINDOW_354,FROM_WINDOW_355,FROM_WINDOW_356,FROM_WINDOW_357,FROM_WINDOW_358,FROM_WINDOW_359,FROM_WINDOW_360,FROM_WINDOW_361,FROM_WINDOW_362,FROM_WINDOW_363,FROM_WINDOW_364,FROM_WINDOW_365,FROM_WINDOW_366,FROM_WINDOW_367,FROM_WINDOW_368,FROM_WINDOW_369,FROM_WINDOW_370,FROM_WINDOW_371,FROM_WINDOW_372,FROM_WINDOW_373,FROM_WINDOW_374,FROM_WINDOW_375,FROM_WINDOW_376,FROM_WINDOW_377,FROM_WINDOW_378,FROM_WINDOW_379,FROM_WINDOW_380,FROM_WINDOW_381,FROM_WINDOW_382,FROM_WINDOW_383,FROM_WINDOW_384,FROM_WINDOW_385,FROM_WINDOW_386,FROM_WINDOW_387,FROM_WINDOW_388,FROM_WINDOW_389,FROM_WINDOW_390,FROM_WINDOW_391,FROM_WINDOW_392,FROM_WINDOW_393,FROM_WINDOW_394,FROM_WINDOW_395,FROM_WINDOW_396,FROM_WINDOW_397,FROM_WINDOW_398,FROM_WINDOW_399,FROM_WINDOW_400,FROM_WINDOW_401,FROM_WINDOW_402,FROM_WINDOW_403,FROM_WINDOW_404,FROM_WINDOW_405,FROM_WINDOW_406,FROM_WINDOW_407,FROM_WINDOW_408,FROM_WINDOW_409,FROM_WINDOW_410,FROM_WINDOW_411,FROM_WINDOW_412,FROM_WINDOW_413,FROM_WINDOW_414,FROM_WINDOW_415,FROM_WINDOW_416,FROM_WINDOW_417,FROM_WINDOW_418,FROM_WINDOW_419,FROM_WINDOW_420,FROM_WINDOW_421,FROM_WINDOW_422,FROM_WINDOW_423,FROM_WINDOW_424,FROM_WINDOW_425,FROM_WINDOW_426,FROM_WINDOW_427,FROM_WINDOW_428,FROM_WINDOW_429,FROM_WINDOW_430,FROM_WINDOW_431,FROM_WINDOW_432,FROM_WINDOW_433,FROM_WINDOW_434,FROM_WINDOW_435,FROM_WINDOW_436,FROM_WINDOW_437,FROM_WINDOW_438,FROM_WINDOW_439,FROM_WINDOW_440,FROM_WINDOW_441,FROM_WINDOW_442,FROM_WINDOW_443,FROM_WINDOW_444,FROM_WINDOW_445,FROM_WINDOW_446,FROM_WINDOW_447,FROM_WINDOW_448,FROM_WINDOW_449,FROM_WINDOW_450,FROM_WINDOW_451,FROM_WINDOW_452,FROM_WINDOW_453,FROM_WINDOW_454,FROM_WINDOW_455,FROM_WINDOW_456,FROM_WINDOW_457,FROM_WINDOW_458,FROM_WINDOW_459,FROM_WINDOW_460,FROM_WINDOW_461,FROM_WINDOW_462,FROM_WINDOW_463,FROM_WINDOW_464,FROM_WINDOW_465,FROM_WINDOW_466,FROM_WINDOW_467,FROM_WINDOW_468,FROM_WINDOW_469,FROM_WINDOW_470,FROM_WINDOW_471,FROM_WINDOW_472,FROM_WINDOW_473,FROM_WINDOW_474,FROM_WINDOW_475,FROM_WINDOW_476,FROM_WINDOW_477,FROM_WINDOW_478,FROM_WINDOW_479,FROM_WINDOW_480,FROM_WINDOW_481,FROM_WINDOW_482,FROM_WINDOW_483,FROM_WINDOW_484,FROM_WINDOW_485,FROM_WINDOW_486,FROM_WINDOW_487,FROM_WINDOW_488,FROM_WINDOW_489,FROM_WINDOW_490,FROM_WINDOW_491,FROM_WINDOW_492,FROM_WINDOW_493,FROM_WINDOW_494,FROM_WINDOW_495,FROM_WINDOW_496,FROM_WINDOW_497,FROM_WINDOW_498,FROM_WINDOW_499,FROM_WINDOW_500,FROM_WINDOW_501,FROM_WINDOW_502,FROM_WINDOW_503,FROM_WINDOW_504,FROM_WINDOW_505,FROM_WINDOW_506,FROM_WINDOW_507,FROM_WINDOW_508,FROM_WINDOW_509,FROM_WINDOW_510,FROM_WINDOW_511,FROM_WINDOW_512,FROM_WINDOW_513,FROM_WINDOW_514,FROM_WINDOW_515,FROM_WINDOW_516,FROM_WINDOW_517,FROM_WINDOW_518,FROM_WINDOW_519,FROM_WINDOW_520,FROM_WINDOW_521,FROM_WINDOW_522,FROM_WINDOW_523,FROM_WINDOW_524,FROM_WINDOW_525,FROM_WINDOW_526,FROM_WINDOW_527,FROM_WINDOW_528,FROM_WINDOW_529,FROM_WINDOW_530,FROM_WINDOW_531,FROM_WINDOW_532,FROM_WINDOW_533,FROM_WINDOW_534,FROM_WINDOW_535,FROM_WINDOW_536,FROM_WINDOW_537,FROM_WINDOW_538,FROM_WINDOW_539,FROM_WINDOW_540,FROM_WINDOW_541,FROM_WINDOW_542,FROM_WINDOW_543,FROM_WINDOW_544,FROM_WINDOW_545,FROM_WINDOW_546,FROM_WINDOW_547,FROM_WINDOW_548,FROM_WINDOW_549,FROM_WINDOW_550,FROM_WINDOW_551,FROM_WINDOW_552,FROM_WINDOW_553,FROM_WINDOW_554,FROM_WINDOW_555,FROM_WINDOW_556,FROM_WINDOW_557,FROM_WINDOW_558,FROM_WINDOW_559,FROM_WINDOW_560,FROM_WINDOW_561,FROM_WINDOW_562,FROM_WINDOW_563,FROM_WINDOW_564,FROM_WINDOW_565,FROM_WINDOW_566,FROM_WINDOW_567,FROM_WINDOW_568,FROM_WINDOW_569,FROM_WINDOW_570,FROM_WINDOW_571,FROM_WINDOW_572,FROM_WINDOW_573,FROM_WINDOW_574,FROM_WINDOW_575,FROM_WINDOW_576,FROM_WINDOW_577,FROM_WINDOW_578,FROM_WINDOW_579,FROM_WINDOW_580,FROM_WINDOW_581,FROM_WINDOW_582,FROM_WINDOW_583,FROM_WINDOW_584,FROM_WINDOW_585,FROM_WINDOW_586,FROM_WINDOW_587,FROM_WINDOW_588,FROM_WINDOW_589,FROM_WINDOW_590,FROM_WINDOW_591,FROM_WINDOW_592,FROM_WINDOW_593,FROM_WINDOW_594,FROM_WINDOW_595,FROM_WINDOW_596,FROM_WINDOW_597,FROM_WINDOW_598,FROM_WINDOW_599,FROM_WINDOW_600,FROM_WINDOW_601,FROM_WINDOW_602,FROM_WINDOW_603,FROM_WINDOW_604,FROM_WINDOW_605,FROM_WINDOW_606,FROM_WINDOW_607,FROM_WINDOW_608,FROM_WINDOW_609,FROM_WINDOW_610,FROM_WINDOW_611,FROM_WINDOW_612,FROM_WINDOW_613,FROM_WINDOW_614,FROM_WINDOW_615,FROM_WINDOW_616,FROM_WINDOW_617,FROM_WINDOW_618,FROM_WINDOW_619,FROM_WINDOW_620,FROM_WINDOW_621,FROM_WINDOW_622,FROM_WINDOW_623,FROM_WINDOW_624,FROM_WINDOW_625,FROM_WINDOW_626,FROM_WINDOW_627,FROM_WINDOW_628,FROM_WINDOW_629,FROM_WINDOW_630,FROM_WINDOW_631,FROM_WINDOW_632,FROM_WINDOW_633,FROM_WINDOW_634,FROM_WINDOW_635,FROM_WINDOW_636,FROM_WINDOW_637,FROM_WINDOW_638,FROM_WINDOW_639,FROM_WINDOW_640,FROM_WINDOW_641,FROM_WINDOW_642,FROM_WINDOW_643,FROM_WINDOW_644,FROM_WINDOW_645,FROM_WINDOW_646,FROM_WINDOW_647,FROM_WINDOW_648,FROM_WINDOW_649,FROM_WINDOW_650,FROM_WINDOW_651,FROM_WINDOW_652,FROM_WINDOW_653,FROM_WINDOW_654,FROM_WINDOW_655,FROM_WINDOW_656,FROM_WINDOW_657,FROM_WINDOW_658,FROM_WINDOW_659,FROM_WINDOW_660,FROM_WINDOW_661,FROM_WINDOW_662,FROM_WINDOW_663,FROM_WINDOW_664,FROM_WINDOW_665,FROM_WINDOW_666,FROM_WINDOW_667,FROM_WINDOW_668,FROM_WINDOW_669,FROM_WINDOW_670,FROM_WINDOW_671,FROM_WINDOW_672,FROM_WINDOW_673,FROM_WINDOW_674,FROM_WINDOW_675,FROM_WINDOW_676,FROM_WINDOW_677,FROM_WINDOW_678,FROM_WINDOW_679,FROM_WINDOW_680,FROM_WINDOW_681,FROM_WINDOW_682,FROM_WINDOW_683,FROM_WINDOW_684,FROM_WINDOW_685,FROM_WINDOW_686,FROM_WINDOW_687,FROM_WINDOW_688,FROM_WINDOW_689,FROM_WINDOW_690,FROM_WINDOW_691,FROM_WINDOW_692,FROM_WINDOW_693,FROM_WINDOW_694,FROM_WINDOW_695,FROM_WINDOW_696,FROM_WINDOW_697,FROM_WINDOW_698,FROM_WINDOW_699,FROM_WINDOW_700,FROM_WINDOW_701,FROM_WINDOW_702,FROM_WINDOW_703,FROM_WINDOW_704,FROM_WINDOW_705,FROM_WINDOW_706,FROM_WINDOW_707,FROM_WINDOW_708,FROM_WINDOW_709,FROM_WINDOW_710,FROM_WINDOW_711,FROM_WINDOW_712,FROM_WINDOW_713,FROM_WINDOW_714,FROM_WINDOW_715,FROM_WINDOW_716,FROM_WINDOW_717,FROM_WINDOW_718,FROM_WINDOW_719,FROM_WINDOW_720,FROM_WINDOW_721,FROM_WINDOW_722,FROM_WINDOW_723,FROM_WINDOW_724,FROM_WINDOW_725,FROM_WINDOW_726,FROM_WINDOW_727,FROM_WINDOW_728,FROM_WINDOW_729,FROM_WINDOW_730,FROM_WINDOW_731,FROM_WINDOW_732,FROM_WINDOW_733,FROM_WINDOW_734,FROM_WINDOW_735,FROM_WINDOW_736,FROM_WINDOW_737,FROM_WINDOW_738,FROM_WINDOW_739,FROM_WINDOW_740,FROM_WINDOW_741,FROM_WINDOW_742,FROM_WINDOW_743,FROM_WINDOW_744,FROM_WINDOW_745,FROM_WINDOW_746,FROM_WINDOW_747,FROM_WINDOW_748,FROM_WINDOW_749,FROM_WINDOW_750,FROM_WINDOW_751,FROM_WINDOW_752,FROM_WINDOW_753,FROM_WINDOW_754,FROM_WINDOW_755,FROM_WINDOW_756,FROM_WINDOW_757,FROM_WINDOW_758,FROM_WINDOW_759,FROM_WINDOW_760,FROM_WINDOW_761,FROM_WINDOW_762,FROM_WINDOW_763,FROM_WINDOW_764,FROM_WINDOW_765,FROM_WINDOW_766,FROM_WINDOW_767,FROM_WINDOW_768,FROM_WINDOW_769,FROM_WINDOW_770,FROM_WINDOW_771,FROM_WINDOW_772,FROM_WINDOW_773,FROM_WINDOW_774,FROM_WINDOW_775,FROM_WINDOW_776,FROM_WINDOW_777,FROM_WINDOW_778,FROM_WINDOW_779,FROM_WINDOW_780,FROM_WINDOW_781,FROM_WINDOW_782,FROM_WINDOW_783,FROM_WINDOW_784,FROM_WINDOW_785,FROM_WINDOW_786,FROM_WINDOW_787,FROM_WINDOW_788,FROM_WINDOW_789,FROM_WINDOW_790,FROM_WINDOW_791,FROM_WINDOW_792,FROM_WINDOW_793,FROM_WINDOW_794,FROM_WINDOW_795,FROM_WINDOW_796,FROM_WINDOW_797,FROM_WINDOW_798,FROM_WINDOW_799,FROM_WINDOW_800,FROM_WINDOW_801,FROM_WINDOW_802,FROM_WINDOW_803,FROM_WINDOW_804,FROM_WINDOW_805,FROM_WINDOW_806,FROM_WINDOW_807,FROM_WINDOW_808,FROM_WINDOW_809,FROM_WINDOW_810,FROM_WINDOW_811,FROM_WINDOW_812,FROM_WINDOW_813,FROM_WINDOW_814,FROM_WINDOW_815,FROM_WINDOW_816,FROM_WINDOW_817,FROM_WINDOW_818,FROM_WINDOW_819,FROM_WINDOW_820,FROM_WINDOW_821,FROM_WINDOW_822,FROM_WINDOW_823,FROM_WINDOW_824,FROM_WINDOW_825,FROM_WINDOW_826,FROM_WINDOW_827,FROM_WINDOW_828,FROM_WINDOW_829,FROM_WINDOW_830,FROM_WINDOW_831,FROM_WINDOW_832,FROM_WINDOW_833,FROM_WINDOW_834,FROM_WINDOW_835,FROM_WINDOW_836,FROM_WINDOW_837,FROM_WINDOW_838,FROM_WINDOW_839,FROM_WINDOW_840,FROM_WINDOW_841,FROM_WINDOW_842,FROM_WINDOW_843,FROM_WINDOW_844,FROM_WINDOW_845,FROM_WINDOW_846,FROM_WINDOW_847,FROM_WINDOW_848,FROM_WINDOW_849,FROM_WINDOW_850,FROM_WINDOW_851,FROM_WINDOW_852,FROM_WINDOW_853,FROM_WINDOW_854,FROM_WINDOW_855,FROM_WINDOW_856,FROM_WINDOW_857,FROM_WINDOW_858,FROM_WINDOW_859,FROM_WINDOW_860,FROM_WINDOW_861,FROM_WINDOW_862,FROM_WINDOW_863,FROM_WINDOW_864,FROM_WINDOW_865,FROM_WINDOW_866,FROM_WINDOW_867,FROM_WINDOW_868,FROM_WINDOW_869,FROM_WINDOW_870,FROM_WINDOW_871,FROM_WINDOW_872,FROM_WINDOW_873,FROM_WINDOW_874,FROM_WINDOW_875,FROM_WINDOW_876,FROM_WINDOW_877,FROM_WINDOW_878,FROM_WINDOW_879,FROM_WINDOW_880,FROM_WINDOW_881,FROM_WINDOW_882,FROM_WINDOW_883,FROM_WINDOW_884,FROM_WINDOW_885,FROM_WINDOW_886,FROM_WINDOW_887,FROM_WINDOW_888,FROM_WINDOW_889,FROM_WINDOW_890,FROM_WINDOW_891,FROM_WINDOW_892,FROM_WINDOW_893,FROM_WINDOW_894,FROM_WINDOW_895,FROM_WINDOW_896,FROM_WINDOW_897,FROM_WINDOW_898,FROM_WINDOW_899,FROM_WINDOW_900,FROM_WINDOW_901,FROM_WINDOW_902,FROM_WINDOW_903,FROM_WINDOW_904,FROM_WINDOW_905,FROM_WINDOW_906,FROM_WINDOW_907,FROM_WINDOW_908,FROM_WINDOW_909,FROM_WINDOW_910,FROM_WINDOW_911,FROM_WINDOW_912,FROM_WINDOW_913,FROM_WINDOW_914,FROM_WINDOW_915,FROM_WINDOW_916,FROM_WINDOW_917,FROM_WINDOW_918,FROM_WINDOW_919,FROM_WINDOW_920,FROM_WINDOW_921,FROM_WINDOW_922,FROM_WINDOW_923,FROM_WINDOW_924,FROM_WINDOW_925,FROM_WINDOW_926,FROM_WINDOW_927,FROM_WINDOW_928,FROM_WINDOW_929,FROM_WINDOW_930,FROM_WINDOW_931,FROM_WINDOW_932,FROM_WINDOW_933,FROM_WINDOW_934,FROM_WINDOW_935,FROM_WINDOW_936,FROM_WINDOW_937,FROM_WINDOW_938,FROM_WINDOW_939,FROM_WINDOW_940,FROM_WINDOW_941,FROM_WINDOW_942,FROM_WINDOW_943,FROM_WINDOW_944,FROM_WINDOW_945,FROM_WINDOW_946,FROM_WINDOW_947,FROM_WINDOW_948,FROM_WINDOW_949,FROM_WINDOW_950,FROM_WINDOW_951,FROM_WINDOW_952,FROM_WINDOW_953,FROM_WINDOW_954,FROM_WINDOW_955,FROM_WINDOW_956,FROM_WINDOW_957,FROM_WINDOW_958,FROM_WINDOW_959,FROM_WINDOW_960,FROM_WINDOW_961,FROM_WINDOW_962,FROM_WINDOW_963,FROM_WINDOW_964,FROM_WINDOW_965,FROM_WINDOW_966,FROM_WINDOW_967,FROM_WINDOW_968,FROM_WINDOW_969,FROM_WINDOW_970,FROM_WINDOW_971,FROM_WINDOW_972,FROM_WINDOW_973,FROM_WINDOW_974,FROM_WINDOW_975,FROM_WINDOW_976,FROM_WINDOW_977,FROM_WINDOW_978,FROM_WINDOW_979,FROM_WINDOW_980,FROM_WINDOW_981,FROM_WINDOW_982,FROM_WINDOW_983,FROM_WINDOW_984,FROM_WINDOW_985,FROM_WINDOW_986,FROM_WINDOW_987,FROM_WINDOW_988,FROM_WINDOW_989,FROM_WINDOW_990,FROM_WINDOW_991,FROM_WINDOW_992,FROM_WINDOW_993,FROM_WINDOW_994,FROM_WINDOW_995,FROM_WINDOW_996,FROM_WINDOW_997,FROM_WINDOW_998,FROM_WINDOW_999,FROM_WINDOW_1000,FROM_WINDOW_1001,FROM_WINDOW_1002,FROM_WINDOW_1003,FROM_WINDOW_1004,FROM_WINDOW_1005,FROM_WINDOW_1006,FROM_WINDOW_1007,FROM_WINDOW_1008,FROM_WINDOW_1009,FROM_WINDOW_1010,FROM_WINDOW_1011,FROM_WINDOW_1012,FROM_WINDOW_1013,FROM_WINDOW_1014,FROM_WINDOW_1015,FROM_WINDOW_1016,FROM_WINDOW_1017,FROM_WINDOW_1018,FROM_WINDOW_1019,FROM_WINDOW_1020,FROM_WINDOW_1021,FROM_WINDOW_1022,FROM_WINDOW_1023: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL MASKED_INPUT_0,MASKED_INPUT_2,MASKED_INPUT_4,MASKED_INPUT_6,MASKED_INPUT_8,MASKED_INPUT_10,MASKED_INPUT_12,MASKED_INPUT_14,MASKED_INPUT_16,MASKED_INPUT_18,MASKED_INPUT_20,MASKED_INPUT_22,MASKED_INPUT_24,MASKED_INPUT_26,MASKED_INPUT_28,MASKED_INPUT_30,MASKED_INPUT_32,MASKED_INPUT_34,MASKED_INPUT_36,MASKED_INPUT_38,MASKED_INPUT_40,MASKED_INPUT_42,MASKED_INPUT_44,MASKED_INPUT_46,MASKED_INPUT_48,MASKED_INPUT_50,MASKED_INPUT_52,MASKED_INPUT_54,MASKED_INPUT_56,MASKED_INPUT_58,MASKED_INPUT_60,MASKED_INPUT_62,MASKED_INPUT_64,MASKED_INPUT_66,MASKED_INPUT_68,MASKED_INPUT_70,MASKED_INPUT_72,MASKED_INPUT_74,MASKED_INPUT_76,MASKED_INPUT_78,MASKED_INPUT_80,MASKED_INPUT_82,MASKED_INPUT_84,MASKED_INPUT_86,MASKED_INPUT_88,MASKED_INPUT_90,MASKED_INPUT_92,MASKED_INPUT_94,MASKED_INPUT_96,MASKED_INPUT_98,MASKED_INPUT_100,MASKED_INPUT_102,MASKED_INPUT_104,MASKED_INPUT_106,MASKED_INPUT_108,MASKED_INPUT_110,MASKED_INPUT_112,MASKED_INPUT_114,MASKED_INPUT_116,MASKED_INPUT_118,MASKED_INPUT_120,MASKED_INPUT_122,MASKED_INPUT_124,MASKED_INPUT_126,MASKED_INPUT_128,MASKED_INPUT_130,MASKED_INPUT_132,MASKED_INPUT_134,MASKED_INPUT_136,MASKED_INPUT_138,MASKED_INPUT_140,MASKED_INPUT_142,MASKED_INPUT_144,MASKED_INPUT_146,MASKED_INPUT_148,MASKED_INPUT_150,MASKED_INPUT_152,MASKED_INPUT_154,MASKED_INPUT_156,MASKED_INPUT_158,MASKED_INPUT_160,MASKED_INPUT_162,MASKED_INPUT_164,MASKED_INPUT_166,MASKED_INPUT_168,MASKED_INPUT_170,MASKED_INPUT_172,MASKED_INPUT_174,MASKED_INPUT_176,MASKED_INPUT_178,MASKED_INPUT_180,MASKED_INPUT_182,MASKED_INPUT_184,MASKED_INPUT_186,MASKED_INPUT_188,MASKED_INPUT_190,MASKED_INPUT_192,MASKED_INPUT_194,MASKED_INPUT_196,MASKED_INPUT_198,MASKED_INPUT_200,MASKED_INPUT_202,MASKED_INPUT_204,MASKED_INPUT_206,MASKED_INPUT_208,MASKED_INPUT_210,MASKED_INPUT_212,MASKED_INPUT_214,MASKED_INPUT_216,MASKED_INPUT_218,MASKED_INPUT_220,MASKED_INPUT_222,MASKED_INPUT_224,MASKED_INPUT_226,MASKED_INPUT_228,MASKED_INPUT_230,MASKED_INPUT_232,MASKED_INPUT_234,MASKED_INPUT_236,MASKED_INPUT_238,MASKED_INPUT_240,MASKED_INPUT_242,MASKED_INPUT_244,MASKED_INPUT_246,MASKED_INPUT_248,MASKED_INPUT_250,MASKED_INPUT_252,MASKED_INPUT_254,MASKED_INPUT_256,MASKED_INPUT_258,MASKED_INPUT_260,MASKED_INPUT_262,MASKED_INPUT_264,MASKED_INPUT_266,MASKED_INPUT_268,MASKED_INPUT_270,MASKED_INPUT_272,MASKED_INPUT_274,MASKED_INPUT_276,MASKED_INPUT_278,MASKED_INPUT_280,MASKED_INPUT_282,MASKED_INPUT_284,MASKED_INPUT_286,MASKED_INPUT_288,MASKED_INPUT_290,MASKED_INPUT_292,MASKED_INPUT_294,MASKED_INPUT_296,MASKED_INPUT_298,MASKED_INPUT_300,MASKED_INPUT_302,MASKED_INPUT_304,MASKED_INPUT_306,MASKED_INPUT_308,MASKED_INPUT_310,MASKED_INPUT_312,MASKED_INPUT_314,MASKED_INPUT_316,MASKED_INPUT_318,MASKED_INPUT_320,MASKED_INPUT_322,MASKED_INPUT_324,MASKED_INPUT_326,MASKED_INPUT_328,MASKED_INPUT_330,MASKED_INPUT_332,MASKED_INPUT_334,MASKED_INPUT_336,MASKED_INPUT_338,MASKED_INPUT_340,MASKED_INPUT_342,MASKED_INPUT_344,MASKED_INPUT_346,MASKED_INPUT_348,MASKED_INPUT_350,MASKED_INPUT_352,MASKED_INPUT_354,MASKED_INPUT_356,MASKED_INPUT_358,MASKED_INPUT_360,MASKED_INPUT_362,MASKED_INPUT_364,MASKED_INPUT_366,MASKED_INPUT_368,MASKED_INPUT_370,MASKED_INPUT_372,MASKED_INPUT_374,MASKED_INPUT_376,MASKED_INPUT_378,MASKED_INPUT_380,MASKED_INPUT_382,MASKED_INPUT_384,MASKED_INPUT_386,MASKED_INPUT_388,MASKED_INPUT_390,MASKED_INPUT_392,MASKED_INPUT_394,MASKED_INPUT_396,MASKED_INPUT_398,MASKED_INPUT_400,MASKED_INPUT_402,MASKED_INPUT_404,MASKED_INPUT_406,MASKED_INPUT_408,MASKED_INPUT_410,MASKED_INPUT_412,MASKED_INPUT_414,MASKED_INPUT_416,MASKED_INPUT_418,MASKED_INPUT_420,MASKED_INPUT_422,MASKED_INPUT_424,MASKED_INPUT_426,MASKED_INPUT_428,MASKED_INPUT_430,MASKED_INPUT_432,MASKED_INPUT_434,MASKED_INPUT_436,MASKED_INPUT_438,MASKED_INPUT_440,MASKED_INPUT_442,MASKED_INPUT_444,MASKED_INPUT_446,MASKED_INPUT_448,MASKED_INPUT_450,MASKED_INPUT_452,MASKED_INPUT_454,MASKED_INPUT_456,MASKED_INPUT_458,MASKED_INPUT_460,MASKED_INPUT_462,MASKED_INPUT_464,MASKED_INPUT_466,MASKED_INPUT_468,MASKED_INPUT_470,MASKED_INPUT_472,MASKED_INPUT_474,MASKED_INPUT_476,MASKED_INPUT_478,MASKED_INPUT_480,MASKED_INPUT_482,MASKED_INPUT_484,MASKED_INPUT_486,MASKED_INPUT_488,MASKED_INPUT_490,MASKED_INPUT_492,MASKED_INPUT_494,MASKED_INPUT_496,MASKED_INPUT_498,MASKED_INPUT_500,MASKED_INPUT_502,MASKED_INPUT_504,MASKED_INPUT_506,MASKED_INPUT_508,MASKED_INPUT_510,MASKED_INPUT_512,MASKED_INPUT_514,MASKED_INPUT_516,MASKED_INPUT_518,MASKED_INPUT_520,MASKED_INPUT_522,MASKED_INPUT_524,MASKED_INPUT_526,MASKED_INPUT_528,MASKED_INPUT_530,MASKED_INPUT_532,MASKED_INPUT_534,MASKED_INPUT_536,MASKED_INPUT_538,MASKED_INPUT_540,MASKED_INPUT_542,MASKED_INPUT_544,MASKED_INPUT_546,MASKED_INPUT_548,MASKED_INPUT_550,MASKED_INPUT_552,MASKED_INPUT_554,MASKED_INPUT_556,MASKED_INPUT_558,MASKED_INPUT_560,MASKED_INPUT_562,MASKED_INPUT_564,MASKED_INPUT_566,MASKED_INPUT_568,MASKED_INPUT_570,MASKED_INPUT_572,MASKED_INPUT_574,MASKED_INPUT_576,MASKED_INPUT_578,MASKED_INPUT_580,MASKED_INPUT_582,MASKED_INPUT_584,MASKED_INPUT_586,MASKED_INPUT_588,MASKED_INPUT_590,MASKED_INPUT_592,MASKED_INPUT_594,MASKED_INPUT_596,MASKED_INPUT_598,MASKED_INPUT_600,MASKED_INPUT_602,MASKED_INPUT_604,MASKED_INPUT_606,MASKED_INPUT_608,MASKED_INPUT_610,MASKED_INPUT_612,MASKED_INPUT_614,MASKED_INPUT_616,MASKED_INPUT_618,MASKED_INPUT_620,MASKED_INPUT_622,MASKED_INPUT_624,MASKED_INPUT_626,MASKED_INPUT_628,MASKED_INPUT_630,MASKED_INPUT_632,MASKED_INPUT_634,MASKED_INPUT_636,MASKED_INPUT_638,MASKED_INPUT_640,MASKED_INPUT_642,MASKED_INPUT_644,MASKED_INPUT_646,MASKED_INPUT_648,MASKED_INPUT_650,MASKED_INPUT_652,MASKED_INPUT_654,MASKED_INPUT_656,MASKED_INPUT_658,MASKED_INPUT_660,MASKED_INPUT_662,MASKED_INPUT_664,MASKED_INPUT_666,MASKED_INPUT_668,MASKED_INPUT_670,MASKED_INPUT_672,MASKED_INPUT_674,MASKED_INPUT_676,MASKED_INPUT_678,MASKED_INPUT_680,MASKED_INPUT_682,MASKED_INPUT_684,MASKED_INPUT_686,MASKED_INPUT_688,MASKED_INPUT_690,MASKED_INPUT_692,MASKED_INPUT_694,MASKED_INPUT_696,MASKED_INPUT_698,MASKED_INPUT_700,MASKED_INPUT_702,MASKED_INPUT_704,MASKED_INPUT_706,MASKED_INPUT_708,MASKED_INPUT_710,MASKED_INPUT_712,MASKED_INPUT_714,MASKED_INPUT_716,MASKED_INPUT_718,MASKED_INPUT_720,MASKED_INPUT_722,MASKED_INPUT_724,MASKED_INPUT_726,MASKED_INPUT_728,MASKED_INPUT_730,MASKED_INPUT_732,MASKED_INPUT_734,MASKED_INPUT_736,MASKED_INPUT_738,MASKED_INPUT_740,MASKED_INPUT_742,MASKED_INPUT_744,MASKED_INPUT_746,MASKED_INPUT_748,MASKED_INPUT_750,MASKED_INPUT_752,MASKED_INPUT_754,MASKED_INPUT_756,MASKED_INPUT_758,MASKED_INPUT_760,MASKED_INPUT_762,MASKED_INPUT_764,MASKED_INPUT_766,MASKED_INPUT_768,MASKED_INPUT_770,MASKED_INPUT_772,MASKED_INPUT_774,MASKED_INPUT_776,MASKED_INPUT_778,MASKED_INPUT_780,MASKED_INPUT_782,MASKED_INPUT_784,MASKED_INPUT_786,MASKED_INPUT_788,MASKED_INPUT_790,MASKED_INPUT_792,MASKED_INPUT_794,MASKED_INPUT_796,MASKED_INPUT_798,MASKED_INPUT_800,MASKED_INPUT_802,MASKED_INPUT_804,MASKED_INPUT_806,MASKED_INPUT_808,MASKED_INPUT_810,MASKED_INPUT_812,MASKED_INPUT_814,MASKED_INPUT_816,MASKED_INPUT_818,MASKED_INPUT_820,MASKED_INPUT_822,MASKED_INPUT_824,MASKED_INPUT_826,MASKED_INPUT_828,MASKED_INPUT_830,MASKED_INPUT_832,MASKED_INPUT_834,MASKED_INPUT_836,MASKED_INPUT_838,MASKED_INPUT_840,MASKED_INPUT_842,MASKED_INPUT_844,MASKED_INPUT_846,MASKED_INPUT_848,MASKED_INPUT_850,MASKED_INPUT_852,MASKED_INPUT_854,MASKED_INPUT_856,MASKED_INPUT_858,MASKED_INPUT_860,MASKED_INPUT_862,MASKED_INPUT_864,MASKED_INPUT_866,MASKED_INPUT_868,MASKED_INPUT_870,MASKED_INPUT_872,MASKED_INPUT_874,MASKED_INPUT_876,MASKED_INPUT_878,MASKED_INPUT_880,MASKED_INPUT_882,MASKED_INPUT_884,MASKED_INPUT_886,MASKED_INPUT_888,MASKED_INPUT_890,MASKED_INPUT_892,MASKED_INPUT_894,MASKED_INPUT_896,MASKED_INPUT_898,MASKED_INPUT_900,MASKED_INPUT_902,MASKED_INPUT_904,MASKED_INPUT_906,MASKED_INPUT_908,MASKED_INPUT_910,MASKED_INPUT_912,MASKED_INPUT_914,MASKED_INPUT_916,MASKED_INPUT_918,MASKED_INPUT_920,MASKED_INPUT_922,MASKED_INPUT_924,MASKED_INPUT_926,MASKED_INPUT_928,MASKED_INPUT_930,MASKED_INPUT_932,MASKED_INPUT_934,MASKED_INPUT_936,MASKED_INPUT_938,MASKED_INPUT_940,MASKED_INPUT_942,MASKED_INPUT_944,MASKED_INPUT_946,MASKED_INPUT_948,MASKED_INPUT_950,MASKED_INPUT_952,MASKED_INPUT_954,MASKED_INPUT_956,MASKED_INPUT_958,MASKED_INPUT_960,MASKED_INPUT_962,MASKED_INPUT_964,MASKED_INPUT_966,MASKED_INPUT_968,MASKED_INPUT_970,MASKED_INPUT_972,MASKED_INPUT_974,MASKED_INPUT_976,MASKED_INPUT_978,MASKED_INPUT_980,MASKED_INPUT_982,MASKED_INPUT_984,MASKED_INPUT_986,MASKED_INPUT_988,MASKED_INPUT_990,MASKED_INPUT_992,MASKED_INPUT_994,MASKED_INPUT_996,MASKED_INPUT_998,MASKED_INPUT_1000,MASKED_INPUT_1002,MASKED_INPUT_1004,MASKED_INPUT_1006,MASKED_INPUT_1008,MASKED_INPUT_1010,MASKED_INPUT_1012,MASKED_INPUT_1014,MASKED_INPUT_1016,MASKED_INPUT_1018,MASKED_INPUT_1020,MASKED_INPUT_1022: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_DATAPATHS_0,FROM_DATAPATHS_1,FROM_DATAPATHS_2,FROM_DATAPATHS_3,FROM_DATAPATHS_4,FROM_DATAPATHS_5,FROM_DATAPATHS_6,FROM_DATAPATHS_7,FROM_DATAPATHS_8,FROM_DATAPATHS_9,FROM_DATAPATHS_10,FROM_DATAPATHS_11,FROM_DATAPATHS_12,FROM_DATAPATHS_13,FROM_DATAPATHS_14,FROM_DATAPATHS_15,FROM_DATAPATHS_16,FROM_DATAPATHS_17,FROM_DATAPATHS_18,FROM_DATAPATHS_19,FROM_DATAPATHS_20,FROM_DATAPATHS_21,FROM_DATAPATHS_22,FROM_DATAPATHS_23,FROM_DATAPATHS_24,FROM_DATAPATHS_25,FROM_DATAPATHS_26,FROM_DATAPATHS_27,FROM_DATAPATHS_28,FROM_DATAPATHS_29,FROM_DATAPATHS_30,FROM_DATAPATHS_31,FROM_DATAPATHS_32,FROM_DATAPATHS_33,FROM_DATAPATHS_34,FROM_DATAPATHS_35,FROM_DATAPATHS_36,FROM_DATAPATHS_37,FROM_DATAPATHS_38,FROM_DATAPATHS_39,FROM_DATAPATHS_40,FROM_DATAPATHS_41,FROM_DATAPATHS_42,FROM_DATAPATHS_43,FROM_DATAPATHS_44,FROM_DATAPATHS_45,FROM_DATAPATHS_46,FROM_DATAPATHS_47,FROM_DATAPATHS_48,FROM_DATAPATHS_49,FROM_DATAPATHS_50,FROM_DATAPATHS_51,FROM_DATAPATHS_52,FROM_DATAPATHS_53,FROM_DATAPATHS_54,FROM_DATAPATHS_55,FROM_DATAPATHS_56,FROM_DATAPATHS_57,FROM_DATAPATHS_58,FROM_DATAPATHS_59,FROM_DATAPATHS_60,FROM_DATAPATHS_61,FROM_DATAPATHS_62,FROM_DATAPATHS_63,FROM_DATAPATHS_64,FROM_DATAPATHS_65,FROM_DATAPATHS_66,FROM_DATAPATHS_67,FROM_DATAPATHS_68,FROM_DATAPATHS_69,FROM_DATAPATHS_70,FROM_DATAPATHS_71,FROM_DATAPATHS_72,FROM_DATAPATHS_73,FROM_DATAPATHS_74,FROM_DATAPATHS_75,FROM_DATAPATHS_76,FROM_DATAPATHS_77,FROM_DATAPATHS_78,FROM_DATAPATHS_79,FROM_DATAPATHS_80,FROM_DATAPATHS_81,FROM_DATAPATHS_82,FROM_DATAPATHS_83,FROM_DATAPATHS_84,FROM_DATAPATHS_85,FROM_DATAPATHS_86,FROM_DATAPATHS_87,FROM_DATAPATHS_88,FROM_DATAPATHS_89,FROM_DATAPATHS_90,FROM_DATAPATHS_91,FROM_DATAPATHS_92,FROM_DATAPATHS_93,FROM_DATAPATHS_94,FROM_DATAPATHS_95,FROM_DATAPATHS_96,FROM_DATAPATHS_97,FROM_DATAPATHS_98,FROM_DATAPATHS_99,FROM_DATAPATHS_100,FROM_DATAPATHS_101,FROM_DATAPATHS_102,FROM_DATAPATHS_103,FROM_DATAPATHS_104,FROM_DATAPATHS_105,FROM_DATAPATHS_106,FROM_DATAPATHS_107,FROM_DATAPATHS_108,FROM_DATAPATHS_109,FROM_DATAPATHS_110,FROM_DATAPATHS_111,FROM_DATAPATHS_112,FROM_DATAPATHS_113,FROM_DATAPATHS_114,FROM_DATAPATHS_115,FROM_DATAPATHS_116,FROM_DATAPATHS_117,FROM_DATAPATHS_118,FROM_DATAPATHS_119,FROM_DATAPATHS_120,FROM_DATAPATHS_121,FROM_DATAPATHS_122,FROM_DATAPATHS_123,FROM_DATAPATHS_124,FROM_DATAPATHS_125,FROM_DATAPATHS_126,FROM_DATAPATHS_127,FROM_DATAPATHS_128,FROM_DATAPATHS_129,FROM_DATAPATHS_130,FROM_DATAPATHS_131,FROM_DATAPATHS_132,FROM_DATAPATHS_133,FROM_DATAPATHS_134,FROM_DATAPATHS_135,FROM_DATAPATHS_136,FROM_DATAPATHS_137,FROM_DATAPATHS_138,FROM_DATAPATHS_139,FROM_DATAPATHS_140,FROM_DATAPATHS_141,FROM_DATAPATHS_142,FROM_DATAPATHS_143,FROM_DATAPATHS_144,FROM_DATAPATHS_145,FROM_DATAPATHS_146,FROM_DATAPATHS_147,FROM_DATAPATHS_148,FROM_DATAPATHS_149,FROM_DATAPATHS_150,FROM_DATAPATHS_151,FROM_DATAPATHS_152,FROM_DATAPATHS_153,FROM_DATAPATHS_154,FROM_DATAPATHS_155,FROM_DATAPATHS_156,FROM_DATAPATHS_157,FROM_DATAPATHS_158,FROM_DATAPATHS_159,FROM_DATAPATHS_160,FROM_DATAPATHS_161,FROM_DATAPATHS_162,FROM_DATAPATHS_163,FROM_DATAPATHS_164,FROM_DATAPATHS_165,FROM_DATAPATHS_166,FROM_DATAPATHS_167,FROM_DATAPATHS_168,FROM_DATAPATHS_169,FROM_DATAPATHS_170,FROM_DATAPATHS_171,FROM_DATAPATHS_172,FROM_DATAPATHS_173,FROM_DATAPATHS_174,FROM_DATAPATHS_175,FROM_DATAPATHS_176,FROM_DATAPATHS_177,FROM_DATAPATHS_178,FROM_DATAPATHS_179,FROM_DATAPATHS_180,FROM_DATAPATHS_181,FROM_DATAPATHS_182,FROM_DATAPATHS_183,FROM_DATAPATHS_184,FROM_DATAPATHS_185,FROM_DATAPATHS_186,FROM_DATAPATHS_187,FROM_DATAPATHS_188,FROM_DATAPATHS_189,FROM_DATAPATHS_190,FROM_DATAPATHS_191,FROM_DATAPATHS_192,FROM_DATAPATHS_193,FROM_DATAPATHS_194,FROM_DATAPATHS_195,FROM_DATAPATHS_196,FROM_DATAPATHS_197,FROM_DATAPATHS_198,FROM_DATAPATHS_199,FROM_DATAPATHS_200,FROM_DATAPATHS_201,FROM_DATAPATHS_202,FROM_DATAPATHS_203,FROM_DATAPATHS_204,FROM_DATAPATHS_205,FROM_DATAPATHS_206,FROM_DATAPATHS_207,FROM_DATAPATHS_208,FROM_DATAPATHS_209,FROM_DATAPATHS_210,FROM_DATAPATHS_211,FROM_DATAPATHS_212,FROM_DATAPATHS_213,FROM_DATAPATHS_214,FROM_DATAPATHS_215,FROM_DATAPATHS_216,FROM_DATAPATHS_217,FROM_DATAPATHS_218,FROM_DATAPATHS_219,FROM_DATAPATHS_220,FROM_DATAPATHS_221,FROM_DATAPATHS_222,FROM_DATAPATHS_223,FROM_DATAPATHS_224,FROM_DATAPATHS_225,FROM_DATAPATHS_226,FROM_DATAPATHS_227,FROM_DATAPATHS_228,FROM_DATAPATHS_229,FROM_DATAPATHS_230,FROM_DATAPATHS_231,FROM_DATAPATHS_232,FROM_DATAPATHS_233,FROM_DATAPATHS_234,FROM_DATAPATHS_235,FROM_DATAPATHS_236,FROM_DATAPATHS_237,FROM_DATAPATHS_238,FROM_DATAPATHS_239,FROM_DATAPATHS_240,FROM_DATAPATHS_241,FROM_DATAPATHS_242,FROM_DATAPATHS_243,FROM_DATAPATHS_244,FROM_DATAPATHS_245,FROM_DATAPATHS_246,FROM_DATAPATHS_247,FROM_DATAPATHS_248,FROM_DATAPATHS_249,FROM_DATAPATHS_250,FROM_DATAPATHS_251,FROM_DATAPATHS_252,FROM_DATAPATHS_253,FROM_DATAPATHS_254,FROM_DATAPATHS_255,FROM_DATAPATHS_256,FROM_DATAPATHS_257,FROM_DATAPATHS_258,FROM_DATAPATHS_259,FROM_DATAPATHS_260,FROM_DATAPATHS_261,FROM_DATAPATHS_262,FROM_DATAPATHS_263,FROM_DATAPATHS_264,FROM_DATAPATHS_265,FROM_DATAPATHS_266,FROM_DATAPATHS_267,FROM_DATAPATHS_268,FROM_DATAPATHS_269,FROM_DATAPATHS_270,FROM_DATAPATHS_271,FROM_DATAPATHS_272,FROM_DATAPATHS_273,FROM_DATAPATHS_274,FROM_DATAPATHS_275,FROM_DATAPATHS_276,FROM_DATAPATHS_277,FROM_DATAPATHS_278,FROM_DATAPATHS_279,FROM_DATAPATHS_280,FROM_DATAPATHS_281,FROM_DATAPATHS_282,FROM_DATAPATHS_283,FROM_DATAPATHS_284,FROM_DATAPATHS_285,FROM_DATAPATHS_286,FROM_DATAPATHS_287,FROM_DATAPATHS_288,FROM_DATAPATHS_289,FROM_DATAPATHS_290,FROM_DATAPATHS_291,FROM_DATAPATHS_292,FROM_DATAPATHS_293,FROM_DATAPATHS_294,FROM_DATAPATHS_295,FROM_DATAPATHS_296,FROM_DATAPATHS_297,FROM_DATAPATHS_298,FROM_DATAPATHS_299,FROM_DATAPATHS_300,FROM_DATAPATHS_301,FROM_DATAPATHS_302,FROM_DATAPATHS_303,FROM_DATAPATHS_304,FROM_DATAPATHS_305,FROM_DATAPATHS_306,FROM_DATAPATHS_307,FROM_DATAPATHS_308,FROM_DATAPATHS_309,FROM_DATAPATHS_310,FROM_DATAPATHS_311,FROM_DATAPATHS_312,FROM_DATAPATHS_313,FROM_DATAPATHS_314,FROM_DATAPATHS_315,FROM_DATAPATHS_316,FROM_DATAPATHS_317,FROM_DATAPATHS_318,FROM_DATAPATHS_319,FROM_DATAPATHS_320,FROM_DATAPATHS_321,FROM_DATAPATHS_322,FROM_DATAPATHS_323,FROM_DATAPATHS_324,FROM_DATAPATHS_325,FROM_DATAPATHS_326,FROM_DATAPATHS_327,FROM_DATAPATHS_328,FROM_DATAPATHS_329,FROM_DATAPATHS_330,FROM_DATAPATHS_331,FROM_DATAPATHS_332,FROM_DATAPATHS_333,FROM_DATAPATHS_334,FROM_DATAPATHS_335,FROM_DATAPATHS_336,FROM_DATAPATHS_337,FROM_DATAPATHS_338,FROM_DATAPATHS_339,FROM_DATAPATHS_340,FROM_DATAPATHS_341,FROM_DATAPATHS_342,FROM_DATAPATHS_343,FROM_DATAPATHS_344,FROM_DATAPATHS_345,FROM_DATAPATHS_346,FROM_DATAPATHS_347,FROM_DATAPATHS_348,FROM_DATAPATHS_349,FROM_DATAPATHS_350,FROM_DATAPATHS_351,FROM_DATAPATHS_352,FROM_DATAPATHS_353,FROM_DATAPATHS_354,FROM_DATAPATHS_355,FROM_DATAPATHS_356,FROM_DATAPATHS_357,FROM_DATAPATHS_358,FROM_DATAPATHS_359,FROM_DATAPATHS_360,FROM_DATAPATHS_361,FROM_DATAPATHS_362,FROM_DATAPATHS_363,FROM_DATAPATHS_364,FROM_DATAPATHS_365,FROM_DATAPATHS_366,FROM_DATAPATHS_367,FROM_DATAPATHS_368,FROM_DATAPATHS_369,FROM_DATAPATHS_370,FROM_DATAPATHS_371,FROM_DATAPATHS_372,FROM_DATAPATHS_373,FROM_DATAPATHS_374,FROM_DATAPATHS_375,FROM_DATAPATHS_376,FROM_DATAPATHS_377,FROM_DATAPATHS_378,FROM_DATAPATHS_379,FROM_DATAPATHS_380,FROM_DATAPATHS_381,FROM_DATAPATHS_382,FROM_DATAPATHS_383,FROM_DATAPATHS_384,FROM_DATAPATHS_385,FROM_DATAPATHS_386,FROM_DATAPATHS_387,FROM_DATAPATHS_388,FROM_DATAPATHS_389,FROM_DATAPATHS_390,FROM_DATAPATHS_391,FROM_DATAPATHS_392,FROM_DATAPATHS_393,FROM_DATAPATHS_394,FROM_DATAPATHS_395,FROM_DATAPATHS_396,FROM_DATAPATHS_397,FROM_DATAPATHS_398,FROM_DATAPATHS_399,FROM_DATAPATHS_400,FROM_DATAPATHS_401,FROM_DATAPATHS_402,FROM_DATAPATHS_403,FROM_DATAPATHS_404,FROM_DATAPATHS_405,FROM_DATAPATHS_406,FROM_DATAPATHS_407,FROM_DATAPATHS_408,FROM_DATAPATHS_409,FROM_DATAPATHS_410,FROM_DATAPATHS_411,FROM_DATAPATHS_412,FROM_DATAPATHS_413,FROM_DATAPATHS_414,FROM_DATAPATHS_415,FROM_DATAPATHS_416,FROM_DATAPATHS_417,FROM_DATAPATHS_418,FROM_DATAPATHS_419,FROM_DATAPATHS_420,FROM_DATAPATHS_421,FROM_DATAPATHS_422,FROM_DATAPATHS_423,FROM_DATAPATHS_424,FROM_DATAPATHS_425,FROM_DATAPATHS_426,FROM_DATAPATHS_427,FROM_DATAPATHS_428,FROM_DATAPATHS_429,FROM_DATAPATHS_430,FROM_DATAPATHS_431,FROM_DATAPATHS_432,FROM_DATAPATHS_433,FROM_DATAPATHS_434,FROM_DATAPATHS_435,FROM_DATAPATHS_436,FROM_DATAPATHS_437,FROM_DATAPATHS_438,FROM_DATAPATHS_439,FROM_DATAPATHS_440,FROM_DATAPATHS_441,FROM_DATAPATHS_442,FROM_DATAPATHS_443,FROM_DATAPATHS_444,FROM_DATAPATHS_445,FROM_DATAPATHS_446,FROM_DATAPATHS_447,FROM_DATAPATHS_448,FROM_DATAPATHS_449,FROM_DATAPATHS_450,FROM_DATAPATHS_451,FROM_DATAPATHS_452,FROM_DATAPATHS_453,FROM_DATAPATHS_454,FROM_DATAPATHS_455,FROM_DATAPATHS_456,FROM_DATAPATHS_457,FROM_DATAPATHS_458,FROM_DATAPATHS_459,FROM_DATAPATHS_460,FROM_DATAPATHS_461,FROM_DATAPATHS_462,FROM_DATAPATHS_463,FROM_DATAPATHS_464,FROM_DATAPATHS_465,FROM_DATAPATHS_466,FROM_DATAPATHS_467,FROM_DATAPATHS_468,FROM_DATAPATHS_469,FROM_DATAPATHS_470,FROM_DATAPATHS_471,FROM_DATAPATHS_472,FROM_DATAPATHS_473,FROM_DATAPATHS_474,FROM_DATAPATHS_475,FROM_DATAPATHS_476,FROM_DATAPATHS_477,FROM_DATAPATHS_478,FROM_DATAPATHS_479,FROM_DATAPATHS_480,FROM_DATAPATHS_481,FROM_DATAPATHS_482,FROM_DATAPATHS_483,FROM_DATAPATHS_484,FROM_DATAPATHS_485,FROM_DATAPATHS_486,FROM_DATAPATHS_487,FROM_DATAPATHS_488,FROM_DATAPATHS_489,FROM_DATAPATHS_490,FROM_DATAPATHS_491,FROM_DATAPATHS_492,FROM_DATAPATHS_493,FROM_DATAPATHS_494,FROM_DATAPATHS_495,FROM_DATAPATHS_496,FROM_DATAPATHS_497,FROM_DATAPATHS_498,FROM_DATAPATHS_499,FROM_DATAPATHS_500,FROM_DATAPATHS_501,FROM_DATAPATHS_502,FROM_DATAPATHS_503,FROM_DATAPATHS_504,FROM_DATAPATHS_505,FROM_DATAPATHS_506,FROM_DATAPATHS_507,FROM_DATAPATHS_508,FROM_DATAPATHS_509,FROM_DATAPATHS_510,FROM_DATAPATHS_511,FROM_DATAPATHS_512,FROM_DATAPATHS_513,FROM_DATAPATHS_514,FROM_DATAPATHS_515,FROM_DATAPATHS_516,FROM_DATAPATHS_517,FROM_DATAPATHS_518,FROM_DATAPATHS_519,FROM_DATAPATHS_520,FROM_DATAPATHS_521,FROM_DATAPATHS_522,FROM_DATAPATHS_523,FROM_DATAPATHS_524,FROM_DATAPATHS_525,FROM_DATAPATHS_526,FROM_DATAPATHS_527,FROM_DATAPATHS_528,FROM_DATAPATHS_529,FROM_DATAPATHS_530,FROM_DATAPATHS_531,FROM_DATAPATHS_532,FROM_DATAPATHS_533,FROM_DATAPATHS_534,FROM_DATAPATHS_535,FROM_DATAPATHS_536,FROM_DATAPATHS_537,FROM_DATAPATHS_538,FROM_DATAPATHS_539,FROM_DATAPATHS_540,FROM_DATAPATHS_541,FROM_DATAPATHS_542,FROM_DATAPATHS_543,FROM_DATAPATHS_544,FROM_DATAPATHS_545,FROM_DATAPATHS_546,FROM_DATAPATHS_547,FROM_DATAPATHS_548,FROM_DATAPATHS_549,FROM_DATAPATHS_550,FROM_DATAPATHS_551,FROM_DATAPATHS_552,FROM_DATAPATHS_553,FROM_DATAPATHS_554,FROM_DATAPATHS_555,FROM_DATAPATHS_556,FROM_DATAPATHS_557,FROM_DATAPATHS_558,FROM_DATAPATHS_559,FROM_DATAPATHS_560,FROM_DATAPATHS_561,FROM_DATAPATHS_562,FROM_DATAPATHS_563,FROM_DATAPATHS_564,FROM_DATAPATHS_565,FROM_DATAPATHS_566,FROM_DATAPATHS_567,FROM_DATAPATHS_568,FROM_DATAPATHS_569,FROM_DATAPATHS_570,FROM_DATAPATHS_571,FROM_DATAPATHS_572,FROM_DATAPATHS_573,FROM_DATAPATHS_574,FROM_DATAPATHS_575,FROM_DATAPATHS_576,FROM_DATAPATHS_577,FROM_DATAPATHS_578,FROM_DATAPATHS_579,FROM_DATAPATHS_580,FROM_DATAPATHS_581,FROM_DATAPATHS_582,FROM_DATAPATHS_583,FROM_DATAPATHS_584,FROM_DATAPATHS_585,FROM_DATAPATHS_586,FROM_DATAPATHS_587,FROM_DATAPATHS_588,FROM_DATAPATHS_589,FROM_DATAPATHS_590,FROM_DATAPATHS_591,FROM_DATAPATHS_592,FROM_DATAPATHS_593,FROM_DATAPATHS_594,FROM_DATAPATHS_595,FROM_DATAPATHS_596,FROM_DATAPATHS_597,FROM_DATAPATHS_598,FROM_DATAPATHS_599,FROM_DATAPATHS_600,FROM_DATAPATHS_601,FROM_DATAPATHS_602,FROM_DATAPATHS_603,FROM_DATAPATHS_604,FROM_DATAPATHS_605,FROM_DATAPATHS_606,FROM_DATAPATHS_607,FROM_DATAPATHS_608,FROM_DATAPATHS_609,FROM_DATAPATHS_610,FROM_DATAPATHS_611,FROM_DATAPATHS_612,FROM_DATAPATHS_613,FROM_DATAPATHS_614,FROM_DATAPATHS_615,FROM_DATAPATHS_616,FROM_DATAPATHS_617,FROM_DATAPATHS_618,FROM_DATAPATHS_619,FROM_DATAPATHS_620,FROM_DATAPATHS_621,FROM_DATAPATHS_622,FROM_DATAPATHS_623,FROM_DATAPATHS_624,FROM_DATAPATHS_625,FROM_DATAPATHS_626,FROM_DATAPATHS_627,FROM_DATAPATHS_628,FROM_DATAPATHS_629,FROM_DATAPATHS_630,FROM_DATAPATHS_631,FROM_DATAPATHS_632,FROM_DATAPATHS_633,FROM_DATAPATHS_634,FROM_DATAPATHS_635,FROM_DATAPATHS_636,FROM_DATAPATHS_637,FROM_DATAPATHS_638,FROM_DATAPATHS_639,FROM_DATAPATHS_640,FROM_DATAPATHS_641,FROM_DATAPATHS_642,FROM_DATAPATHS_643,FROM_DATAPATHS_644,FROM_DATAPATHS_645,FROM_DATAPATHS_646,FROM_DATAPATHS_647,FROM_DATAPATHS_648,FROM_DATAPATHS_649,FROM_DATAPATHS_650,FROM_DATAPATHS_651,FROM_DATAPATHS_652,FROM_DATAPATHS_653,FROM_DATAPATHS_654,FROM_DATAPATHS_655,FROM_DATAPATHS_656,FROM_DATAPATHS_657,FROM_DATAPATHS_658,FROM_DATAPATHS_659,FROM_DATAPATHS_660,FROM_DATAPATHS_661,FROM_DATAPATHS_662,FROM_DATAPATHS_663,FROM_DATAPATHS_664,FROM_DATAPATHS_665,FROM_DATAPATHS_666,FROM_DATAPATHS_667,FROM_DATAPATHS_668,FROM_DATAPATHS_669,FROM_DATAPATHS_670,FROM_DATAPATHS_671,FROM_DATAPATHS_672,FROM_DATAPATHS_673,FROM_DATAPATHS_674,FROM_DATAPATHS_675,FROM_DATAPATHS_676,FROM_DATAPATHS_677,FROM_DATAPATHS_678,FROM_DATAPATHS_679,FROM_DATAPATHS_680,FROM_DATAPATHS_681,FROM_DATAPATHS_682,FROM_DATAPATHS_683,FROM_DATAPATHS_684,FROM_DATAPATHS_685,FROM_DATAPATHS_686,FROM_DATAPATHS_687,FROM_DATAPATHS_688,FROM_DATAPATHS_689,FROM_DATAPATHS_690,FROM_DATAPATHS_691,FROM_DATAPATHS_692,FROM_DATAPATHS_693,FROM_DATAPATHS_694,FROM_DATAPATHS_695,FROM_DATAPATHS_696,FROM_DATAPATHS_697,FROM_DATAPATHS_698,FROM_DATAPATHS_699,FROM_DATAPATHS_700,FROM_DATAPATHS_701,FROM_DATAPATHS_702,FROM_DATAPATHS_703,FROM_DATAPATHS_704,FROM_DATAPATHS_705,FROM_DATAPATHS_706,FROM_DATAPATHS_707,FROM_DATAPATHS_708,FROM_DATAPATHS_709,FROM_DATAPATHS_710,FROM_DATAPATHS_711,FROM_DATAPATHS_712,FROM_DATAPATHS_713,FROM_DATAPATHS_714,FROM_DATAPATHS_715,FROM_DATAPATHS_716,FROM_DATAPATHS_717,FROM_DATAPATHS_718,FROM_DATAPATHS_719,FROM_DATAPATHS_720,FROM_DATAPATHS_721,FROM_DATAPATHS_722,FROM_DATAPATHS_723,FROM_DATAPATHS_724,FROM_DATAPATHS_725,FROM_DATAPATHS_726,FROM_DATAPATHS_727,FROM_DATAPATHS_728,FROM_DATAPATHS_729,FROM_DATAPATHS_730,FROM_DATAPATHS_731,FROM_DATAPATHS_732,FROM_DATAPATHS_733,FROM_DATAPATHS_734,FROM_DATAPATHS_735,FROM_DATAPATHS_736,FROM_DATAPATHS_737,FROM_DATAPATHS_738,FROM_DATAPATHS_739,FROM_DATAPATHS_740,FROM_DATAPATHS_741,FROM_DATAPATHS_742,FROM_DATAPATHS_743,FROM_DATAPATHS_744,FROM_DATAPATHS_745,FROM_DATAPATHS_746,FROM_DATAPATHS_747,FROM_DATAPATHS_748,FROM_DATAPATHS_749,FROM_DATAPATHS_750,FROM_DATAPATHS_751,FROM_DATAPATHS_752,FROM_DATAPATHS_753,FROM_DATAPATHS_754,FROM_DATAPATHS_755,FROM_DATAPATHS_756,FROM_DATAPATHS_757,FROM_DATAPATHS_758,FROM_DATAPATHS_759,FROM_DATAPATHS_760,FROM_DATAPATHS_761,FROM_DATAPATHS_762,FROM_DATAPATHS_763,FROM_DATAPATHS_764,FROM_DATAPATHS_765,FROM_DATAPATHS_766,FROM_DATAPATHS_767,FROM_DATAPATHS_768,FROM_DATAPATHS_769,FROM_DATAPATHS_770,FROM_DATAPATHS_771,FROM_DATAPATHS_772,FROM_DATAPATHS_773,FROM_DATAPATHS_774,FROM_DATAPATHS_775,FROM_DATAPATHS_776,FROM_DATAPATHS_777,FROM_DATAPATHS_778,FROM_DATAPATHS_779,FROM_DATAPATHS_780,FROM_DATAPATHS_781,FROM_DATAPATHS_782,FROM_DATAPATHS_783,FROM_DATAPATHS_784,FROM_DATAPATHS_785,FROM_DATAPATHS_786,FROM_DATAPATHS_787,FROM_DATAPATHS_788,FROM_DATAPATHS_789,FROM_DATAPATHS_790,FROM_DATAPATHS_791,FROM_DATAPATHS_792,FROM_DATAPATHS_793,FROM_DATAPATHS_794,FROM_DATAPATHS_795,FROM_DATAPATHS_796,FROM_DATAPATHS_797,FROM_DATAPATHS_798,FROM_DATAPATHS_799,FROM_DATAPATHS_800,FROM_DATAPATHS_801,FROM_DATAPATHS_802,FROM_DATAPATHS_803,FROM_DATAPATHS_804,FROM_DATAPATHS_805,FROM_DATAPATHS_806,FROM_DATAPATHS_807,FROM_DATAPATHS_808,FROM_DATAPATHS_809,FROM_DATAPATHS_810,FROM_DATAPATHS_811,FROM_DATAPATHS_812,FROM_DATAPATHS_813,FROM_DATAPATHS_814,FROM_DATAPATHS_815,FROM_DATAPATHS_816,FROM_DATAPATHS_817,FROM_DATAPATHS_818,FROM_DATAPATHS_819,FROM_DATAPATHS_820,FROM_DATAPATHS_821,FROM_DATAPATHS_822,FROM_DATAPATHS_823,FROM_DATAPATHS_824,FROM_DATAPATHS_825,FROM_DATAPATHS_826,FROM_DATAPATHS_827,FROM_DATAPATHS_828,FROM_DATAPATHS_829,FROM_DATAPATHS_830,FROM_DATAPATHS_831,FROM_DATAPATHS_832,FROM_DATAPATHS_833,FROM_DATAPATHS_834,FROM_DATAPATHS_835,FROM_DATAPATHS_836,FROM_DATAPATHS_837,FROM_DATAPATHS_838,FROM_DATAPATHS_839,FROM_DATAPATHS_840,FROM_DATAPATHS_841,FROM_DATAPATHS_842,FROM_DATAPATHS_843,FROM_DATAPATHS_844,FROM_DATAPATHS_845,FROM_DATAPATHS_846,FROM_DATAPATHS_847,FROM_DATAPATHS_848,FROM_DATAPATHS_849,FROM_DATAPATHS_850,FROM_DATAPATHS_851,FROM_DATAPATHS_852,FROM_DATAPATHS_853,FROM_DATAPATHS_854,FROM_DATAPATHS_855,FROM_DATAPATHS_856,FROM_DATAPATHS_857,FROM_DATAPATHS_858,FROM_DATAPATHS_859,FROM_DATAPATHS_860,FROM_DATAPATHS_861,FROM_DATAPATHS_862,FROM_DATAPATHS_863,FROM_DATAPATHS_864,FROM_DATAPATHS_865,FROM_DATAPATHS_866,FROM_DATAPATHS_867,FROM_DATAPATHS_868,FROM_DATAPATHS_869,FROM_DATAPATHS_870,FROM_DATAPATHS_871,FROM_DATAPATHS_872,FROM_DATAPATHS_873,FROM_DATAPATHS_874,FROM_DATAPATHS_875,FROM_DATAPATHS_876,FROM_DATAPATHS_877,FROM_DATAPATHS_878,FROM_DATAPATHS_879,FROM_DATAPATHS_880,FROM_DATAPATHS_881,FROM_DATAPATHS_882,FROM_DATAPATHS_883,FROM_DATAPATHS_884,FROM_DATAPATHS_885,FROM_DATAPATHS_886,FROM_DATAPATHS_887,FROM_DATAPATHS_888,FROM_DATAPATHS_889,FROM_DATAPATHS_890,FROM_DATAPATHS_891,FROM_DATAPATHS_892,FROM_DATAPATHS_893,FROM_DATAPATHS_894,FROM_DATAPATHS_895,FROM_DATAPATHS_896,FROM_DATAPATHS_897,FROM_DATAPATHS_898,FROM_DATAPATHS_899,FROM_DATAPATHS_900,FROM_DATAPATHS_901,FROM_DATAPATHS_902,FROM_DATAPATHS_903,FROM_DATAPATHS_904,FROM_DATAPATHS_905,FROM_DATAPATHS_906,FROM_DATAPATHS_907,FROM_DATAPATHS_908,FROM_DATAPATHS_909,FROM_DATAPATHS_910,FROM_DATAPATHS_911,FROM_DATAPATHS_912,FROM_DATAPATHS_913,FROM_DATAPATHS_914,FROM_DATAPATHS_915,FROM_DATAPATHS_916,FROM_DATAPATHS_917,FROM_DATAPATHS_918,FROM_DATAPATHS_919,FROM_DATAPATHS_920,FROM_DATAPATHS_921,FROM_DATAPATHS_922,FROM_DATAPATHS_923,FROM_DATAPATHS_924,FROM_DATAPATHS_925,FROM_DATAPATHS_926,FROM_DATAPATHS_927,FROM_DATAPATHS_928,FROM_DATAPATHS_929,FROM_DATAPATHS_930,FROM_DATAPATHS_931,FROM_DATAPATHS_932,FROM_DATAPATHS_933,FROM_DATAPATHS_934,FROM_DATAPATHS_935,FROM_DATAPATHS_936,FROM_DATAPATHS_937,FROM_DATAPATHS_938,FROM_DATAPATHS_939,FROM_DATAPATHS_940,FROM_DATAPATHS_941,FROM_DATAPATHS_942,FROM_DATAPATHS_943,FROM_DATAPATHS_944,FROM_DATAPATHS_945,FROM_DATAPATHS_946,FROM_DATAPATHS_947,FROM_DATAPATHS_948,FROM_DATAPATHS_949,FROM_DATAPATHS_950,FROM_DATAPATHS_951,FROM_DATAPATHS_952,FROM_DATAPATHS_953,FROM_DATAPATHS_954,FROM_DATAPATHS_955,FROM_DATAPATHS_956,FROM_DATAPATHS_957,FROM_DATAPATHS_958,FROM_DATAPATHS_959,FROM_DATAPATHS_960,FROM_DATAPATHS_961,FROM_DATAPATHS_962,FROM_DATAPATHS_963,FROM_DATAPATHS_964,FROM_DATAPATHS_965,FROM_DATAPATHS_966,FROM_DATAPATHS_967,FROM_DATAPATHS_968,FROM_DATAPATHS_969,FROM_DATAPATHS_970,FROM_DATAPATHS_971,FROM_DATAPATHS_972,FROM_DATAPATHS_973,FROM_DATAPATHS_974,FROM_DATAPATHS_975,FROM_DATAPATHS_976,FROM_DATAPATHS_977,FROM_DATAPATHS_978,FROM_DATAPATHS_979,FROM_DATAPATHS_980,FROM_DATAPATHS_981,FROM_DATAPATHS_982,FROM_DATAPATHS_983,FROM_DATAPATHS_984,FROM_DATAPATHS_985,FROM_DATAPATHS_986,FROM_DATAPATHS_987,FROM_DATAPATHS_988,FROM_DATAPATHS_989,FROM_DATAPATHS_990,FROM_DATAPATHS_991,FROM_DATAPATHS_992,FROM_DATAPATHS_993,FROM_DATAPATHS_994,FROM_DATAPATHS_995,FROM_DATAPATHS_996,FROM_DATAPATHS_997,FROM_DATAPATHS_998,FROM_DATAPATHS_999,FROM_DATAPATHS_1000,FROM_DATAPATHS_1001,FROM_DATAPATHS_1002,FROM_DATAPATHS_1003,FROM_DATAPATHS_1004,FROM_DATAPATHS_1005,FROM_DATAPATHS_1006,FROM_DATAPATHS_1007,FROM_DATAPATHS_1008,FROM_DATAPATHS_1009,FROM_DATAPATHS_1010,FROM_DATAPATHS_1011,FROM_DATAPATHS_1012,FROM_DATAPATHS_1013,FROM_DATAPATHS_1014,FROM_DATAPATHS_1015,FROM_DATAPATHS_1016,FROM_DATAPATHS_1017,FROM_DATAPATHS_1018,FROM_DATAPATHS_1019,FROM_DATAPATHS_1020,FROM_DATAPATHS_1021,FROM_DATAPATHS_1022,FROM_DATAPATHS_1023: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_CONTROL_UNITS_0,FROM_CONTROL_UNITS_1,FROM_CONTROL_UNITS_2,FROM_CONTROL_UNITS_3,FROM_CONTROL_UNITS_4,FROM_CONTROL_UNITS_5,FROM_CONTROL_UNITS_6,FROM_CONTROL_UNITS_7,FROM_CONTROL_UNITS_8,FROM_CONTROL_UNITS_9,FROM_CONTROL_UNITS_10,FROM_CONTROL_UNITS_11,FROM_CONTROL_UNITS_12,FROM_CONTROL_UNITS_13,FROM_CONTROL_UNITS_14,FROM_CONTROL_UNITS_15,FROM_CONTROL_UNITS_16,FROM_CONTROL_UNITS_17,FROM_CONTROL_UNITS_18,FROM_CONTROL_UNITS_19,FROM_CONTROL_UNITS_20,FROM_CONTROL_UNITS_21,FROM_CONTROL_UNITS_22,FROM_CONTROL_UNITS_23,FROM_CONTROL_UNITS_24,FROM_CONTROL_UNITS_25,FROM_CONTROL_UNITS_26,FROM_CONTROL_UNITS_27,FROM_CONTROL_UNITS_28,FROM_CONTROL_UNITS_29,FROM_CONTROL_UNITS_30,FROM_CONTROL_UNITS_31,FROM_CONTROL_UNITS_32,FROM_CONTROL_UNITS_33,FROM_CONTROL_UNITS_34,FROM_CONTROL_UNITS_35,FROM_CONTROL_UNITS_36,FROM_CONTROL_UNITS_37,FROM_CONTROL_UNITS_38,FROM_CONTROL_UNITS_39,FROM_CONTROL_UNITS_40,FROM_CONTROL_UNITS_41,FROM_CONTROL_UNITS_42,FROM_CONTROL_UNITS_43,FROM_CONTROL_UNITS_44,FROM_CONTROL_UNITS_45,FROM_CONTROL_UNITS_46,FROM_CONTROL_UNITS_47,FROM_CONTROL_UNITS_48,FROM_CONTROL_UNITS_49,FROM_CONTROL_UNITS_50,FROM_CONTROL_UNITS_51,FROM_CONTROL_UNITS_52,FROM_CONTROL_UNITS_53,FROM_CONTROL_UNITS_54,FROM_CONTROL_UNITS_55,FROM_CONTROL_UNITS_56,FROM_CONTROL_UNITS_57,FROM_CONTROL_UNITS_58,FROM_CONTROL_UNITS_59,FROM_CONTROL_UNITS_60,FROM_CONTROL_UNITS_61,FROM_CONTROL_UNITS_62,FROM_CONTROL_UNITS_63,FROM_CONTROL_UNITS_64,FROM_CONTROL_UNITS_65,FROM_CONTROL_UNITS_66,FROM_CONTROL_UNITS_67,FROM_CONTROL_UNITS_68,FROM_CONTROL_UNITS_69,FROM_CONTROL_UNITS_70,FROM_CONTROL_UNITS_71,FROM_CONTROL_UNITS_72,FROM_CONTROL_UNITS_73,FROM_CONTROL_UNITS_74,FROM_CONTROL_UNITS_75,FROM_CONTROL_UNITS_76,FROM_CONTROL_UNITS_77,FROM_CONTROL_UNITS_78,FROM_CONTROL_UNITS_79,FROM_CONTROL_UNITS_80,FROM_CONTROL_UNITS_81,FROM_CONTROL_UNITS_82,FROM_CONTROL_UNITS_83,FROM_CONTROL_UNITS_84,FROM_CONTROL_UNITS_85,FROM_CONTROL_UNITS_86,FROM_CONTROL_UNITS_87,FROM_CONTROL_UNITS_88,FROM_CONTROL_UNITS_89,FROM_CONTROL_UNITS_90,FROM_CONTROL_UNITS_91,FROM_CONTROL_UNITS_92,FROM_CONTROL_UNITS_93,FROM_CONTROL_UNITS_94,FROM_CONTROL_UNITS_95,FROM_CONTROL_UNITS_96,FROM_CONTROL_UNITS_97,FROM_CONTROL_UNITS_98,FROM_CONTROL_UNITS_99,FROM_CONTROL_UNITS_100,FROM_CONTROL_UNITS_101,FROM_CONTROL_UNITS_102,FROM_CONTROL_UNITS_103,FROM_CONTROL_UNITS_104,FROM_CONTROL_UNITS_105,FROM_CONTROL_UNITS_106,FROM_CONTROL_UNITS_107,FROM_CONTROL_UNITS_108,FROM_CONTROL_UNITS_109,FROM_CONTROL_UNITS_110,FROM_CONTROL_UNITS_111,FROM_CONTROL_UNITS_112,FROM_CONTROL_UNITS_113,FROM_CONTROL_UNITS_114,FROM_CONTROL_UNITS_115,FROM_CONTROL_UNITS_116,FROM_CONTROL_UNITS_117,FROM_CONTROL_UNITS_118,FROM_CONTROL_UNITS_119,FROM_CONTROL_UNITS_120,FROM_CONTROL_UNITS_121,FROM_CONTROL_UNITS_122,FROM_CONTROL_UNITS_123,FROM_CONTROL_UNITS_124,FROM_CONTROL_UNITS_125,FROM_CONTROL_UNITS_126,FROM_CONTROL_UNITS_127,FROM_CONTROL_UNITS_128,FROM_CONTROL_UNITS_129,FROM_CONTROL_UNITS_130,FROM_CONTROL_UNITS_131,FROM_CONTROL_UNITS_132,FROM_CONTROL_UNITS_133,FROM_CONTROL_UNITS_134,FROM_CONTROL_UNITS_135,FROM_CONTROL_UNITS_136,FROM_CONTROL_UNITS_137,FROM_CONTROL_UNITS_138,FROM_CONTROL_UNITS_139,FROM_CONTROL_UNITS_140,FROM_CONTROL_UNITS_141,FROM_CONTROL_UNITS_142,FROM_CONTROL_UNITS_143,FROM_CONTROL_UNITS_144,FROM_CONTROL_UNITS_145,FROM_CONTROL_UNITS_146,FROM_CONTROL_UNITS_147,FROM_CONTROL_UNITS_148,FROM_CONTROL_UNITS_149,FROM_CONTROL_UNITS_150,FROM_CONTROL_UNITS_151,FROM_CONTROL_UNITS_152,FROM_CONTROL_UNITS_153,FROM_CONTROL_UNITS_154,FROM_CONTROL_UNITS_155,FROM_CONTROL_UNITS_156,FROM_CONTROL_UNITS_157,FROM_CONTROL_UNITS_158,FROM_CONTROL_UNITS_159,FROM_CONTROL_UNITS_160,FROM_CONTROL_UNITS_161,FROM_CONTROL_UNITS_162,FROM_CONTROL_UNITS_163,FROM_CONTROL_UNITS_164,FROM_CONTROL_UNITS_165,FROM_CONTROL_UNITS_166,FROM_CONTROL_UNITS_167,FROM_CONTROL_UNITS_168,FROM_CONTROL_UNITS_169,FROM_CONTROL_UNITS_170,FROM_CONTROL_UNITS_171,FROM_CONTROL_UNITS_172,FROM_CONTROL_UNITS_173,FROM_CONTROL_UNITS_174,FROM_CONTROL_UNITS_175,FROM_CONTROL_UNITS_176,FROM_CONTROL_UNITS_177,FROM_CONTROL_UNITS_178,FROM_CONTROL_UNITS_179,FROM_CONTROL_UNITS_180,FROM_CONTROL_UNITS_181,FROM_CONTROL_UNITS_182,FROM_CONTROL_UNITS_183,FROM_CONTROL_UNITS_184,FROM_CONTROL_UNITS_185,FROM_CONTROL_UNITS_186,FROM_CONTROL_UNITS_187,FROM_CONTROL_UNITS_188,FROM_CONTROL_UNITS_189,FROM_CONTROL_UNITS_190,FROM_CONTROL_UNITS_191,FROM_CONTROL_UNITS_192,FROM_CONTROL_UNITS_193,FROM_CONTROL_UNITS_194,FROM_CONTROL_UNITS_195,FROM_CONTROL_UNITS_196,FROM_CONTROL_UNITS_197,FROM_CONTROL_UNITS_198,FROM_CONTROL_UNITS_199,FROM_CONTROL_UNITS_200,FROM_CONTROL_UNITS_201,FROM_CONTROL_UNITS_202,FROM_CONTROL_UNITS_203,FROM_CONTROL_UNITS_204,FROM_CONTROL_UNITS_205,FROM_CONTROL_UNITS_206,FROM_CONTROL_UNITS_207,FROM_CONTROL_UNITS_208,FROM_CONTROL_UNITS_209,FROM_CONTROL_UNITS_210,FROM_CONTROL_UNITS_211,FROM_CONTROL_UNITS_212,FROM_CONTROL_UNITS_213,FROM_CONTROL_UNITS_214,FROM_CONTROL_UNITS_215,FROM_CONTROL_UNITS_216,FROM_CONTROL_UNITS_217,FROM_CONTROL_UNITS_218,FROM_CONTROL_UNITS_219,FROM_CONTROL_UNITS_220,FROM_CONTROL_UNITS_221,FROM_CONTROL_UNITS_222,FROM_CONTROL_UNITS_223,FROM_CONTROL_UNITS_224,FROM_CONTROL_UNITS_225,FROM_CONTROL_UNITS_226,FROM_CONTROL_UNITS_227,FROM_CONTROL_UNITS_228,FROM_CONTROL_UNITS_229,FROM_CONTROL_UNITS_230,FROM_CONTROL_UNITS_231,FROM_CONTROL_UNITS_232,FROM_CONTROL_UNITS_233,FROM_CONTROL_UNITS_234,FROM_CONTROL_UNITS_235,FROM_CONTROL_UNITS_236,FROM_CONTROL_UNITS_237,FROM_CONTROL_UNITS_238,FROM_CONTROL_UNITS_239,FROM_CONTROL_UNITS_240,FROM_CONTROL_UNITS_241,FROM_CONTROL_UNITS_242,FROM_CONTROL_UNITS_243,FROM_CONTROL_UNITS_244,FROM_CONTROL_UNITS_245,FROM_CONTROL_UNITS_246,FROM_CONTROL_UNITS_247,FROM_CONTROL_UNITS_248,FROM_CONTROL_UNITS_249,FROM_CONTROL_UNITS_250,FROM_CONTROL_UNITS_251,FROM_CONTROL_UNITS_252,FROM_CONTROL_UNITS_253,FROM_CONTROL_UNITS_254,FROM_CONTROL_UNITS_255,FROM_CONTROL_UNITS_256,FROM_CONTROL_UNITS_257,FROM_CONTROL_UNITS_258,FROM_CONTROL_UNITS_259,FROM_CONTROL_UNITS_260,FROM_CONTROL_UNITS_261,FROM_CONTROL_UNITS_262,FROM_CONTROL_UNITS_263,FROM_CONTROL_UNITS_264,FROM_CONTROL_UNITS_265,FROM_CONTROL_UNITS_266,FROM_CONTROL_UNITS_267,FROM_CONTROL_UNITS_268,FROM_CONTROL_UNITS_269,FROM_CONTROL_UNITS_270,FROM_CONTROL_UNITS_271,FROM_CONTROL_UNITS_272,FROM_CONTROL_UNITS_273,FROM_CONTROL_UNITS_274,FROM_CONTROL_UNITS_275,FROM_CONTROL_UNITS_276,FROM_CONTROL_UNITS_277,FROM_CONTROL_UNITS_278,FROM_CONTROL_UNITS_279,FROM_CONTROL_UNITS_280,FROM_CONTROL_UNITS_281,FROM_CONTROL_UNITS_282,FROM_CONTROL_UNITS_283,FROM_CONTROL_UNITS_284,FROM_CONTROL_UNITS_285,FROM_CONTROL_UNITS_286,FROM_CONTROL_UNITS_287,FROM_CONTROL_UNITS_288,FROM_CONTROL_UNITS_289,FROM_CONTROL_UNITS_290,FROM_CONTROL_UNITS_291,FROM_CONTROL_UNITS_292,FROM_CONTROL_UNITS_293,FROM_CONTROL_UNITS_294,FROM_CONTROL_UNITS_295,FROM_CONTROL_UNITS_296,FROM_CONTROL_UNITS_297,FROM_CONTROL_UNITS_298,FROM_CONTROL_UNITS_299,FROM_CONTROL_UNITS_300,FROM_CONTROL_UNITS_301,FROM_CONTROL_UNITS_302,FROM_CONTROL_UNITS_303,FROM_CONTROL_UNITS_304,FROM_CONTROL_UNITS_305,FROM_CONTROL_UNITS_306,FROM_CONTROL_UNITS_307,FROM_CONTROL_UNITS_308,FROM_CONTROL_UNITS_309,FROM_CONTROL_UNITS_310,FROM_CONTROL_UNITS_311,FROM_CONTROL_UNITS_312,FROM_CONTROL_UNITS_313,FROM_CONTROL_UNITS_314,FROM_CONTROL_UNITS_315,FROM_CONTROL_UNITS_316,FROM_CONTROL_UNITS_317,FROM_CONTROL_UNITS_318,FROM_CONTROL_UNITS_319,FROM_CONTROL_UNITS_320,FROM_CONTROL_UNITS_321,FROM_CONTROL_UNITS_322,FROM_CONTROL_UNITS_323,FROM_CONTROL_UNITS_324,FROM_CONTROL_UNITS_325,FROM_CONTROL_UNITS_326,FROM_CONTROL_UNITS_327,FROM_CONTROL_UNITS_328,FROM_CONTROL_UNITS_329,FROM_CONTROL_UNITS_330,FROM_CONTROL_UNITS_331,FROM_CONTROL_UNITS_332,FROM_CONTROL_UNITS_333,FROM_CONTROL_UNITS_334,FROM_CONTROL_UNITS_335,FROM_CONTROL_UNITS_336,FROM_CONTROL_UNITS_337,FROM_CONTROL_UNITS_338,FROM_CONTROL_UNITS_339,FROM_CONTROL_UNITS_340,FROM_CONTROL_UNITS_341,FROM_CONTROL_UNITS_342,FROM_CONTROL_UNITS_343,FROM_CONTROL_UNITS_344,FROM_CONTROL_UNITS_345,FROM_CONTROL_UNITS_346,FROM_CONTROL_UNITS_347,FROM_CONTROL_UNITS_348,FROM_CONTROL_UNITS_349,FROM_CONTROL_UNITS_350,FROM_CONTROL_UNITS_351,FROM_CONTROL_UNITS_352,FROM_CONTROL_UNITS_353,FROM_CONTROL_UNITS_354,FROM_CONTROL_UNITS_355,FROM_CONTROL_UNITS_356,FROM_CONTROL_UNITS_357,FROM_CONTROL_UNITS_358,FROM_CONTROL_UNITS_359,FROM_CONTROL_UNITS_360,FROM_CONTROL_UNITS_361,FROM_CONTROL_UNITS_362,FROM_CONTROL_UNITS_363,FROM_CONTROL_UNITS_364,FROM_CONTROL_UNITS_365,FROM_CONTROL_UNITS_366,FROM_CONTROL_UNITS_367,FROM_CONTROL_UNITS_368,FROM_CONTROL_UNITS_369,FROM_CONTROL_UNITS_370,FROM_CONTROL_UNITS_371,FROM_CONTROL_UNITS_372,FROM_CONTROL_UNITS_373,FROM_CONTROL_UNITS_374,FROM_CONTROL_UNITS_375,FROM_CONTROL_UNITS_376,FROM_CONTROL_UNITS_377,FROM_CONTROL_UNITS_378,FROM_CONTROL_UNITS_379,FROM_CONTROL_UNITS_380,FROM_CONTROL_UNITS_381,FROM_CONTROL_UNITS_382,FROM_CONTROL_UNITS_383,FROM_CONTROL_UNITS_384,FROM_CONTROL_UNITS_385,FROM_CONTROL_UNITS_386,FROM_CONTROL_UNITS_387,FROM_CONTROL_UNITS_388,FROM_CONTROL_UNITS_389,FROM_CONTROL_UNITS_390,FROM_CONTROL_UNITS_391,FROM_CONTROL_UNITS_392,FROM_CONTROL_UNITS_393,FROM_CONTROL_UNITS_394,FROM_CONTROL_UNITS_395,FROM_CONTROL_UNITS_396,FROM_CONTROL_UNITS_397,FROM_CONTROL_UNITS_398,FROM_CONTROL_UNITS_399,FROM_CONTROL_UNITS_400,FROM_CONTROL_UNITS_401,FROM_CONTROL_UNITS_402,FROM_CONTROL_UNITS_403,FROM_CONTROL_UNITS_404,FROM_CONTROL_UNITS_405,FROM_CONTROL_UNITS_406,FROM_CONTROL_UNITS_407,FROM_CONTROL_UNITS_408,FROM_CONTROL_UNITS_409,FROM_CONTROL_UNITS_410,FROM_CONTROL_UNITS_411,FROM_CONTROL_UNITS_412,FROM_CONTROL_UNITS_413,FROM_CONTROL_UNITS_414,FROM_CONTROL_UNITS_415,FROM_CONTROL_UNITS_416,FROM_CONTROL_UNITS_417,FROM_CONTROL_UNITS_418,FROM_CONTROL_UNITS_419,FROM_CONTROL_UNITS_420,FROM_CONTROL_UNITS_421,FROM_CONTROL_UNITS_422,FROM_CONTROL_UNITS_423,FROM_CONTROL_UNITS_424,FROM_CONTROL_UNITS_425,FROM_CONTROL_UNITS_426,FROM_CONTROL_UNITS_427,FROM_CONTROL_UNITS_428,FROM_CONTROL_UNITS_429,FROM_CONTROL_UNITS_430,FROM_CONTROL_UNITS_431,FROM_CONTROL_UNITS_432,FROM_CONTROL_UNITS_433,FROM_CONTROL_UNITS_434,FROM_CONTROL_UNITS_435,FROM_CONTROL_UNITS_436,FROM_CONTROL_UNITS_437,FROM_CONTROL_UNITS_438,FROM_CONTROL_UNITS_439,FROM_CONTROL_UNITS_440,FROM_CONTROL_UNITS_441,FROM_CONTROL_UNITS_442,FROM_CONTROL_UNITS_443,FROM_CONTROL_UNITS_444,FROM_CONTROL_UNITS_445,FROM_CONTROL_UNITS_446,FROM_CONTROL_UNITS_447,FROM_CONTROL_UNITS_448,FROM_CONTROL_UNITS_449,FROM_CONTROL_UNITS_450,FROM_CONTROL_UNITS_451,FROM_CONTROL_UNITS_452,FROM_CONTROL_UNITS_453,FROM_CONTROL_UNITS_454,FROM_CONTROL_UNITS_455,FROM_CONTROL_UNITS_456,FROM_CONTROL_UNITS_457,FROM_CONTROL_UNITS_458,FROM_CONTROL_UNITS_459,FROM_CONTROL_UNITS_460,FROM_CONTROL_UNITS_461,FROM_CONTROL_UNITS_462,FROM_CONTROL_UNITS_463,FROM_CONTROL_UNITS_464,FROM_CONTROL_UNITS_465,FROM_CONTROL_UNITS_466,FROM_CONTROL_UNITS_467,FROM_CONTROL_UNITS_468,FROM_CONTROL_UNITS_469,FROM_CONTROL_UNITS_470,FROM_CONTROL_UNITS_471,FROM_CONTROL_UNITS_472,FROM_CONTROL_UNITS_473,FROM_CONTROL_UNITS_474,FROM_CONTROL_UNITS_475,FROM_CONTROL_UNITS_476,FROM_CONTROL_UNITS_477,FROM_CONTROL_UNITS_478,FROM_CONTROL_UNITS_479,FROM_CONTROL_UNITS_480,FROM_CONTROL_UNITS_481,FROM_CONTROL_UNITS_482,FROM_CONTROL_UNITS_483,FROM_CONTROL_UNITS_484,FROM_CONTROL_UNITS_485,FROM_CONTROL_UNITS_486,FROM_CONTROL_UNITS_487,FROM_CONTROL_UNITS_488,FROM_CONTROL_UNITS_489,FROM_CONTROL_UNITS_490,FROM_CONTROL_UNITS_491,FROM_CONTROL_UNITS_492,FROM_CONTROL_UNITS_493,FROM_CONTROL_UNITS_494,FROM_CONTROL_UNITS_495,FROM_CONTROL_UNITS_496,FROM_CONTROL_UNITS_497,FROM_CONTROL_UNITS_498,FROM_CONTROL_UNITS_499,FROM_CONTROL_UNITS_500,FROM_CONTROL_UNITS_501,FROM_CONTROL_UNITS_502,FROM_CONTROL_UNITS_503,FROM_CONTROL_UNITS_504,FROM_CONTROL_UNITS_505,FROM_CONTROL_UNITS_506,FROM_CONTROL_UNITS_507,FROM_CONTROL_UNITS_508,FROM_CONTROL_UNITS_509,FROM_CONTROL_UNITS_510,FROM_CONTROL_UNITS_511,FROM_CONTROL_UNITS_512,FROM_CONTROL_UNITS_513,FROM_CONTROL_UNITS_514,FROM_CONTROL_UNITS_515,FROM_CONTROL_UNITS_516,FROM_CONTROL_UNITS_517,FROM_CONTROL_UNITS_518,FROM_CONTROL_UNITS_519,FROM_CONTROL_UNITS_520,FROM_CONTROL_UNITS_521,FROM_CONTROL_UNITS_522,FROM_CONTROL_UNITS_523,FROM_CONTROL_UNITS_524,FROM_CONTROL_UNITS_525,FROM_CONTROL_UNITS_526,FROM_CONTROL_UNITS_527,FROM_CONTROL_UNITS_528,FROM_CONTROL_UNITS_529,FROM_CONTROL_UNITS_530,FROM_CONTROL_UNITS_531,FROM_CONTROL_UNITS_532,FROM_CONTROL_UNITS_533,FROM_CONTROL_UNITS_534,FROM_CONTROL_UNITS_535,FROM_CONTROL_UNITS_536,FROM_CONTROL_UNITS_537,FROM_CONTROL_UNITS_538,FROM_CONTROL_UNITS_539,FROM_CONTROL_UNITS_540,FROM_CONTROL_UNITS_541,FROM_CONTROL_UNITS_542,FROM_CONTROL_UNITS_543,FROM_CONTROL_UNITS_544,FROM_CONTROL_UNITS_545,FROM_CONTROL_UNITS_546,FROM_CONTROL_UNITS_547,FROM_CONTROL_UNITS_548,FROM_CONTROL_UNITS_549,FROM_CONTROL_UNITS_550,FROM_CONTROL_UNITS_551,FROM_CONTROL_UNITS_552,FROM_CONTROL_UNITS_553,FROM_CONTROL_UNITS_554,FROM_CONTROL_UNITS_555,FROM_CONTROL_UNITS_556,FROM_CONTROL_UNITS_557,FROM_CONTROL_UNITS_558,FROM_CONTROL_UNITS_559,FROM_CONTROL_UNITS_560,FROM_CONTROL_UNITS_561,FROM_CONTROL_UNITS_562,FROM_CONTROL_UNITS_563,FROM_CONTROL_UNITS_564,FROM_CONTROL_UNITS_565,FROM_CONTROL_UNITS_566,FROM_CONTROL_UNITS_567,FROM_CONTROL_UNITS_568,FROM_CONTROL_UNITS_569,FROM_CONTROL_UNITS_570,FROM_CONTROL_UNITS_571,FROM_CONTROL_UNITS_572,FROM_CONTROL_UNITS_573,FROM_CONTROL_UNITS_574,FROM_CONTROL_UNITS_575,FROM_CONTROL_UNITS_576,FROM_CONTROL_UNITS_577,FROM_CONTROL_UNITS_578,FROM_CONTROL_UNITS_579,FROM_CONTROL_UNITS_580,FROM_CONTROL_UNITS_581,FROM_CONTROL_UNITS_582,FROM_CONTROL_UNITS_583,FROM_CONTROL_UNITS_584,FROM_CONTROL_UNITS_585,FROM_CONTROL_UNITS_586,FROM_CONTROL_UNITS_587,FROM_CONTROL_UNITS_588,FROM_CONTROL_UNITS_589,FROM_CONTROL_UNITS_590,FROM_CONTROL_UNITS_591,FROM_CONTROL_UNITS_592,FROM_CONTROL_UNITS_593,FROM_CONTROL_UNITS_594,FROM_CONTROL_UNITS_595,FROM_CONTROL_UNITS_596,FROM_CONTROL_UNITS_597,FROM_CONTROL_UNITS_598,FROM_CONTROL_UNITS_599,FROM_CONTROL_UNITS_600,FROM_CONTROL_UNITS_601,FROM_CONTROL_UNITS_602,FROM_CONTROL_UNITS_603,FROM_CONTROL_UNITS_604,FROM_CONTROL_UNITS_605,FROM_CONTROL_UNITS_606,FROM_CONTROL_UNITS_607,FROM_CONTROL_UNITS_608,FROM_CONTROL_UNITS_609,FROM_CONTROL_UNITS_610,FROM_CONTROL_UNITS_611,FROM_CONTROL_UNITS_612,FROM_CONTROL_UNITS_613,FROM_CONTROL_UNITS_614,FROM_CONTROL_UNITS_615,FROM_CONTROL_UNITS_616,FROM_CONTROL_UNITS_617,FROM_CONTROL_UNITS_618,FROM_CONTROL_UNITS_619,FROM_CONTROL_UNITS_620,FROM_CONTROL_UNITS_621,FROM_CONTROL_UNITS_622,FROM_CONTROL_UNITS_623,FROM_CONTROL_UNITS_624,FROM_CONTROL_UNITS_625,FROM_CONTROL_UNITS_626,FROM_CONTROL_UNITS_627,FROM_CONTROL_UNITS_628,FROM_CONTROL_UNITS_629,FROM_CONTROL_UNITS_630,FROM_CONTROL_UNITS_631,FROM_CONTROL_UNITS_632,FROM_CONTROL_UNITS_633,FROM_CONTROL_UNITS_634,FROM_CONTROL_UNITS_635,FROM_CONTROL_UNITS_636,FROM_CONTROL_UNITS_637,FROM_CONTROL_UNITS_638,FROM_CONTROL_UNITS_639,FROM_CONTROL_UNITS_640,FROM_CONTROL_UNITS_641,FROM_CONTROL_UNITS_642,FROM_CONTROL_UNITS_643,FROM_CONTROL_UNITS_644,FROM_CONTROL_UNITS_645,FROM_CONTROL_UNITS_646,FROM_CONTROL_UNITS_647,FROM_CONTROL_UNITS_648,FROM_CONTROL_UNITS_649,FROM_CONTROL_UNITS_650,FROM_CONTROL_UNITS_651,FROM_CONTROL_UNITS_652,FROM_CONTROL_UNITS_653,FROM_CONTROL_UNITS_654,FROM_CONTROL_UNITS_655,FROM_CONTROL_UNITS_656,FROM_CONTROL_UNITS_657,FROM_CONTROL_UNITS_658,FROM_CONTROL_UNITS_659,FROM_CONTROL_UNITS_660,FROM_CONTROL_UNITS_661,FROM_CONTROL_UNITS_662,FROM_CONTROL_UNITS_663,FROM_CONTROL_UNITS_664,FROM_CONTROL_UNITS_665,FROM_CONTROL_UNITS_666,FROM_CONTROL_UNITS_667,FROM_CONTROL_UNITS_668,FROM_CONTROL_UNITS_669,FROM_CONTROL_UNITS_670,FROM_CONTROL_UNITS_671,FROM_CONTROL_UNITS_672,FROM_CONTROL_UNITS_673,FROM_CONTROL_UNITS_674,FROM_CONTROL_UNITS_675,FROM_CONTROL_UNITS_676,FROM_CONTROL_UNITS_677,FROM_CONTROL_UNITS_678,FROM_CONTROL_UNITS_679,FROM_CONTROL_UNITS_680,FROM_CONTROL_UNITS_681,FROM_CONTROL_UNITS_682,FROM_CONTROL_UNITS_683,FROM_CONTROL_UNITS_684,FROM_CONTROL_UNITS_685,FROM_CONTROL_UNITS_686,FROM_CONTROL_UNITS_687,FROM_CONTROL_UNITS_688,FROM_CONTROL_UNITS_689,FROM_CONTROL_UNITS_690,FROM_CONTROL_UNITS_691,FROM_CONTROL_UNITS_692,FROM_CONTROL_UNITS_693,FROM_CONTROL_UNITS_694,FROM_CONTROL_UNITS_695,FROM_CONTROL_UNITS_696,FROM_CONTROL_UNITS_697,FROM_CONTROL_UNITS_698,FROM_CONTROL_UNITS_699,FROM_CONTROL_UNITS_700,FROM_CONTROL_UNITS_701,FROM_CONTROL_UNITS_702,FROM_CONTROL_UNITS_703,FROM_CONTROL_UNITS_704,FROM_CONTROL_UNITS_705,FROM_CONTROL_UNITS_706,FROM_CONTROL_UNITS_707,FROM_CONTROL_UNITS_708,FROM_CONTROL_UNITS_709,FROM_CONTROL_UNITS_710,FROM_CONTROL_UNITS_711,FROM_CONTROL_UNITS_712,FROM_CONTROL_UNITS_713,FROM_CONTROL_UNITS_714,FROM_CONTROL_UNITS_715,FROM_CONTROL_UNITS_716,FROM_CONTROL_UNITS_717,FROM_CONTROL_UNITS_718,FROM_CONTROL_UNITS_719,FROM_CONTROL_UNITS_720,FROM_CONTROL_UNITS_721,FROM_CONTROL_UNITS_722,FROM_CONTROL_UNITS_723,FROM_CONTROL_UNITS_724,FROM_CONTROL_UNITS_725,FROM_CONTROL_UNITS_726,FROM_CONTROL_UNITS_727,FROM_CONTROL_UNITS_728,FROM_CONTROL_UNITS_729,FROM_CONTROL_UNITS_730,FROM_CONTROL_UNITS_731,FROM_CONTROL_UNITS_732,FROM_CONTROL_UNITS_733,FROM_CONTROL_UNITS_734,FROM_CONTROL_UNITS_735,FROM_CONTROL_UNITS_736,FROM_CONTROL_UNITS_737,FROM_CONTROL_UNITS_738,FROM_CONTROL_UNITS_739,FROM_CONTROL_UNITS_740,FROM_CONTROL_UNITS_741,FROM_CONTROL_UNITS_742,FROM_CONTROL_UNITS_743,FROM_CONTROL_UNITS_744,FROM_CONTROL_UNITS_745,FROM_CONTROL_UNITS_746,FROM_CONTROL_UNITS_747,FROM_CONTROL_UNITS_748,FROM_CONTROL_UNITS_749,FROM_CONTROL_UNITS_750,FROM_CONTROL_UNITS_751,FROM_CONTROL_UNITS_752,FROM_CONTROL_UNITS_753,FROM_CONTROL_UNITS_754,FROM_CONTROL_UNITS_755,FROM_CONTROL_UNITS_756,FROM_CONTROL_UNITS_757,FROM_CONTROL_UNITS_758,FROM_CONTROL_UNITS_759,FROM_CONTROL_UNITS_760,FROM_CONTROL_UNITS_761,FROM_CONTROL_UNITS_762,FROM_CONTROL_UNITS_763,FROM_CONTROL_UNITS_764,FROM_CONTROL_UNITS_765,FROM_CONTROL_UNITS_766,FROM_CONTROL_UNITS_767,FROM_CONTROL_UNITS_768,FROM_CONTROL_UNITS_769,FROM_CONTROL_UNITS_770,FROM_CONTROL_UNITS_771,FROM_CONTROL_UNITS_772,FROM_CONTROL_UNITS_773,FROM_CONTROL_UNITS_774,FROM_CONTROL_UNITS_775,FROM_CONTROL_UNITS_776,FROM_CONTROL_UNITS_777,FROM_CONTROL_UNITS_778,FROM_CONTROL_UNITS_779,FROM_CONTROL_UNITS_780,FROM_CONTROL_UNITS_781,FROM_CONTROL_UNITS_782,FROM_CONTROL_UNITS_783,FROM_CONTROL_UNITS_784,FROM_CONTROL_UNITS_785,FROM_CONTROL_UNITS_786,FROM_CONTROL_UNITS_787,FROM_CONTROL_UNITS_788,FROM_CONTROL_UNITS_789,FROM_CONTROL_UNITS_790,FROM_CONTROL_UNITS_791,FROM_CONTROL_UNITS_792,FROM_CONTROL_UNITS_793,FROM_CONTROL_UNITS_794,FROM_CONTROL_UNITS_795,FROM_CONTROL_UNITS_796,FROM_CONTROL_UNITS_797,FROM_CONTROL_UNITS_798,FROM_CONTROL_UNITS_799,FROM_CONTROL_UNITS_800,FROM_CONTROL_UNITS_801,FROM_CONTROL_UNITS_802,FROM_CONTROL_UNITS_803,FROM_CONTROL_UNITS_804,FROM_CONTROL_UNITS_805,FROM_CONTROL_UNITS_806,FROM_CONTROL_UNITS_807,FROM_CONTROL_UNITS_808,FROM_CONTROL_UNITS_809,FROM_CONTROL_UNITS_810,FROM_CONTROL_UNITS_811,FROM_CONTROL_UNITS_812,FROM_CONTROL_UNITS_813,FROM_CONTROL_UNITS_814,FROM_CONTROL_UNITS_815,FROM_CONTROL_UNITS_816,FROM_CONTROL_UNITS_817,FROM_CONTROL_UNITS_818,FROM_CONTROL_UNITS_819,FROM_CONTROL_UNITS_820,FROM_CONTROL_UNITS_821,FROM_CONTROL_UNITS_822,FROM_CONTROL_UNITS_823,FROM_CONTROL_UNITS_824,FROM_CONTROL_UNITS_825,FROM_CONTROL_UNITS_826,FROM_CONTROL_UNITS_827,FROM_CONTROL_UNITS_828,FROM_CONTROL_UNITS_829,FROM_CONTROL_UNITS_830,FROM_CONTROL_UNITS_831,FROM_CONTROL_UNITS_832,FROM_CONTROL_UNITS_833,FROM_CONTROL_UNITS_834,FROM_CONTROL_UNITS_835,FROM_CONTROL_UNITS_836,FROM_CONTROL_UNITS_837,FROM_CONTROL_UNITS_838,FROM_CONTROL_UNITS_839,FROM_CONTROL_UNITS_840,FROM_CONTROL_UNITS_841,FROM_CONTROL_UNITS_842,FROM_CONTROL_UNITS_843,FROM_CONTROL_UNITS_844,FROM_CONTROL_UNITS_845,FROM_CONTROL_UNITS_846,FROM_CONTROL_UNITS_847,FROM_CONTROL_UNITS_848,FROM_CONTROL_UNITS_849,FROM_CONTROL_UNITS_850,FROM_CONTROL_UNITS_851,FROM_CONTROL_UNITS_852,FROM_CONTROL_UNITS_853,FROM_CONTROL_UNITS_854,FROM_CONTROL_UNITS_855,FROM_CONTROL_UNITS_856,FROM_CONTROL_UNITS_857,FROM_CONTROL_UNITS_858,FROM_CONTROL_UNITS_859,FROM_CONTROL_UNITS_860,FROM_CONTROL_UNITS_861,FROM_CONTROL_UNITS_862,FROM_CONTROL_UNITS_863,FROM_CONTROL_UNITS_864,FROM_CONTROL_UNITS_865,FROM_CONTROL_UNITS_866,FROM_CONTROL_UNITS_867,FROM_CONTROL_UNITS_868,FROM_CONTROL_UNITS_869,FROM_CONTROL_UNITS_870,FROM_CONTROL_UNITS_871,FROM_CONTROL_UNITS_872,FROM_CONTROL_UNITS_873,FROM_CONTROL_UNITS_874,FROM_CONTROL_UNITS_875,FROM_CONTROL_UNITS_876,FROM_CONTROL_UNITS_877,FROM_CONTROL_UNITS_878,FROM_CONTROL_UNITS_879,FROM_CONTROL_UNITS_880,FROM_CONTROL_UNITS_881,FROM_CONTROL_UNITS_882,FROM_CONTROL_UNITS_883,FROM_CONTROL_UNITS_884,FROM_CONTROL_UNITS_885,FROM_CONTROL_UNITS_886,FROM_CONTROL_UNITS_887,FROM_CONTROL_UNITS_888,FROM_CONTROL_UNITS_889,FROM_CONTROL_UNITS_890,FROM_CONTROL_UNITS_891,FROM_CONTROL_UNITS_892,FROM_CONTROL_UNITS_893,FROM_CONTROL_UNITS_894,FROM_CONTROL_UNITS_895,FROM_CONTROL_UNITS_896,FROM_CONTROL_UNITS_897,FROM_CONTROL_UNITS_898,FROM_CONTROL_UNITS_899,FROM_CONTROL_UNITS_900,FROM_CONTROL_UNITS_901,FROM_CONTROL_UNITS_902,FROM_CONTROL_UNITS_903,FROM_CONTROL_UNITS_904,FROM_CONTROL_UNITS_905,FROM_CONTROL_UNITS_906,FROM_CONTROL_UNITS_907,FROM_CONTROL_UNITS_908,FROM_CONTROL_UNITS_909,FROM_CONTROL_UNITS_910,FROM_CONTROL_UNITS_911,FROM_CONTROL_UNITS_912,FROM_CONTROL_UNITS_913,FROM_CONTROL_UNITS_914,FROM_CONTROL_UNITS_915,FROM_CONTROL_UNITS_916,FROM_CONTROL_UNITS_917,FROM_CONTROL_UNITS_918,FROM_CONTROL_UNITS_919,FROM_CONTROL_UNITS_920,FROM_CONTROL_UNITS_921,FROM_CONTROL_UNITS_922,FROM_CONTROL_UNITS_923,FROM_CONTROL_UNITS_924,FROM_CONTROL_UNITS_925,FROM_CONTROL_UNITS_926,FROM_CONTROL_UNITS_927,FROM_CONTROL_UNITS_928,FROM_CONTROL_UNITS_929,FROM_CONTROL_UNITS_930,FROM_CONTROL_UNITS_931,FROM_CONTROL_UNITS_932,FROM_CONTROL_UNITS_933,FROM_CONTROL_UNITS_934,FROM_CONTROL_UNITS_935,FROM_CONTROL_UNITS_936,FROM_CONTROL_UNITS_937,FROM_CONTROL_UNITS_938,FROM_CONTROL_UNITS_939,FROM_CONTROL_UNITS_940,FROM_CONTROL_UNITS_941,FROM_CONTROL_UNITS_942,FROM_CONTROL_UNITS_943,FROM_CONTROL_UNITS_944,FROM_CONTROL_UNITS_945,FROM_CONTROL_UNITS_946,FROM_CONTROL_UNITS_947,FROM_CONTROL_UNITS_948,FROM_CONTROL_UNITS_949,FROM_CONTROL_UNITS_950,FROM_CONTROL_UNITS_951,FROM_CONTROL_UNITS_952,FROM_CONTROL_UNITS_953,FROM_CONTROL_UNITS_954,FROM_CONTROL_UNITS_955,FROM_CONTROL_UNITS_956,FROM_CONTROL_UNITS_957,FROM_CONTROL_UNITS_958,FROM_CONTROL_UNITS_959,FROM_CONTROL_UNITS_960,FROM_CONTROL_UNITS_961,FROM_CONTROL_UNITS_962,FROM_CONTROL_UNITS_963,FROM_CONTROL_UNITS_964,FROM_CONTROL_UNITS_965,FROM_CONTROL_UNITS_966,FROM_CONTROL_UNITS_967,FROM_CONTROL_UNITS_968,FROM_CONTROL_UNITS_969,FROM_CONTROL_UNITS_970,FROM_CONTROL_UNITS_971,FROM_CONTROL_UNITS_972,FROM_CONTROL_UNITS_973,FROM_CONTROL_UNITS_974,FROM_CONTROL_UNITS_975,FROM_CONTROL_UNITS_976,FROM_CONTROL_UNITS_977,FROM_CONTROL_UNITS_978,FROM_CONTROL_UNITS_979,FROM_CONTROL_UNITS_980,FROM_CONTROL_UNITS_981,FROM_CONTROL_UNITS_982,FROM_CONTROL_UNITS_983,FROM_CONTROL_UNITS_984,FROM_CONTROL_UNITS_985,FROM_CONTROL_UNITS_986,FROM_CONTROL_UNITS_987,FROM_CONTROL_UNITS_988,FROM_CONTROL_UNITS_989,FROM_CONTROL_UNITS_990,FROM_CONTROL_UNITS_991,FROM_CONTROL_UNITS_992,FROM_CONTROL_UNITS_993,FROM_CONTROL_UNITS_994,FROM_CONTROL_UNITS_995,FROM_CONTROL_UNITS_996,FROM_CONTROL_UNITS_997,FROM_CONTROL_UNITS_998,FROM_CONTROL_UNITS_999,FROM_CONTROL_UNITS_1000,FROM_CONTROL_UNITS_1001,FROM_CONTROL_UNITS_1002,FROM_CONTROL_UNITS_1003,FROM_CONTROL_UNITS_1004,FROM_CONTROL_UNITS_1005,FROM_CONTROL_UNITS_1006,FROM_CONTROL_UNITS_1007,FROM_CONTROL_UNITS_1008,FROM_CONTROL_UNITS_1009,FROM_CONTROL_UNITS_1010,FROM_CONTROL_UNITS_1011,FROM_CONTROL_UNITS_1012,FROM_CONTROL_UNITS_1013,FROM_CONTROL_UNITS_1014,FROM_CONTROL_UNITS_1015,FROM_CONTROL_UNITS_1016,FROM_CONTROL_UNITS_1017,FROM_CONTROL_UNITS_1018,FROM_CONTROL_UNITS_1019,FROM_CONTROL_UNITS_1020,FROM_CONTROL_UNITS_1021,FROM_CONTROL_UNITS_1022,FROM_CONTROL_UNITS_1023: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL UNWINDOWED_0,UNWINDOWED_1,UNWINDOWED_2,UNWINDOWED_3,UNWINDOWED_4,UNWINDOWED_5,UNWINDOWED_6,UNWINDOWED_7,UNWINDOWED_8,UNWINDOWED_9,UNWINDOWED_10,UNWINDOWED_11,UNWINDOWED_12,UNWINDOWED_13,UNWINDOWED_14,UNWINDOWED_15,UNWINDOWED_16,UNWINDOWED_17,UNWINDOWED_18,UNWINDOWED_19,UNWINDOWED_20,UNWINDOWED_21,UNWINDOWED_22,UNWINDOWED_23,UNWINDOWED_24,UNWINDOWED_25,UNWINDOWED_26,UNWINDOWED_27,UNWINDOWED_28,UNWINDOWED_29,UNWINDOWED_30,UNWINDOWED_31,UNWINDOWED_32,UNWINDOWED_33,UNWINDOWED_34,UNWINDOWED_35,UNWINDOWED_36,UNWINDOWED_37,UNWINDOWED_38,UNWINDOWED_39,UNWINDOWED_40,UNWINDOWED_41,UNWINDOWED_42,UNWINDOWED_43,UNWINDOWED_44,UNWINDOWED_45,UNWINDOWED_46,UNWINDOWED_47,UNWINDOWED_48,UNWINDOWED_49,UNWINDOWED_50,UNWINDOWED_51,UNWINDOWED_52,UNWINDOWED_53,UNWINDOWED_54,UNWINDOWED_55,UNWINDOWED_56,UNWINDOWED_57,UNWINDOWED_58,UNWINDOWED_59,UNWINDOWED_60,UNWINDOWED_61,UNWINDOWED_62,UNWINDOWED_63,UNWINDOWED_64,UNWINDOWED_65,UNWINDOWED_66,UNWINDOWED_67,UNWINDOWED_68,UNWINDOWED_69,UNWINDOWED_70,UNWINDOWED_71,UNWINDOWED_72,UNWINDOWED_73,UNWINDOWED_74,UNWINDOWED_75,UNWINDOWED_76,UNWINDOWED_77,UNWINDOWED_78,UNWINDOWED_79,UNWINDOWED_80,UNWINDOWED_81,UNWINDOWED_82,UNWINDOWED_83,UNWINDOWED_84,UNWINDOWED_85,UNWINDOWED_86,UNWINDOWED_87,UNWINDOWED_88,UNWINDOWED_89,UNWINDOWED_90,UNWINDOWED_91,UNWINDOWED_92,UNWINDOWED_93,UNWINDOWED_94,UNWINDOWED_95,UNWINDOWED_96,UNWINDOWED_97,UNWINDOWED_98,UNWINDOWED_99,UNWINDOWED_100,UNWINDOWED_101,UNWINDOWED_102,UNWINDOWED_103,UNWINDOWED_104,UNWINDOWED_105,UNWINDOWED_106,UNWINDOWED_107,UNWINDOWED_108,UNWINDOWED_109,UNWINDOWED_110,UNWINDOWED_111,UNWINDOWED_112,UNWINDOWED_113,UNWINDOWED_114,UNWINDOWED_115,UNWINDOWED_116,UNWINDOWED_117,UNWINDOWED_118,UNWINDOWED_119,UNWINDOWED_120,UNWINDOWED_121,UNWINDOWED_122,UNWINDOWED_123,UNWINDOWED_124,UNWINDOWED_125,UNWINDOWED_126,UNWINDOWED_127,UNWINDOWED_128,UNWINDOWED_129,UNWINDOWED_130,UNWINDOWED_131,UNWINDOWED_132,UNWINDOWED_133,UNWINDOWED_134,UNWINDOWED_135,UNWINDOWED_136,UNWINDOWED_137,UNWINDOWED_138,UNWINDOWED_139,UNWINDOWED_140,UNWINDOWED_141,UNWINDOWED_142,UNWINDOWED_143,UNWINDOWED_144,UNWINDOWED_145,UNWINDOWED_146,UNWINDOWED_147,UNWINDOWED_148,UNWINDOWED_149,UNWINDOWED_150,UNWINDOWED_151,UNWINDOWED_152,UNWINDOWED_153,UNWINDOWED_154,UNWINDOWED_155,UNWINDOWED_156,UNWINDOWED_157,UNWINDOWED_158,UNWINDOWED_159,UNWINDOWED_160,UNWINDOWED_161,UNWINDOWED_162,UNWINDOWED_163,UNWINDOWED_164,UNWINDOWED_165,UNWINDOWED_166,UNWINDOWED_167,UNWINDOWED_168,UNWINDOWED_169,UNWINDOWED_170,UNWINDOWED_171,UNWINDOWED_172,UNWINDOWED_173,UNWINDOWED_174,UNWINDOWED_175,UNWINDOWED_176,UNWINDOWED_177,UNWINDOWED_178,UNWINDOWED_179,UNWINDOWED_180,UNWINDOWED_181,UNWINDOWED_182,UNWINDOWED_183,UNWINDOWED_184,UNWINDOWED_185,UNWINDOWED_186,UNWINDOWED_187,UNWINDOWED_188,UNWINDOWED_189,UNWINDOWED_190,UNWINDOWED_191,UNWINDOWED_192,UNWINDOWED_193,UNWINDOWED_194,UNWINDOWED_195,UNWINDOWED_196,UNWINDOWED_197,UNWINDOWED_198,UNWINDOWED_199,UNWINDOWED_200,UNWINDOWED_201,UNWINDOWED_202,UNWINDOWED_203,UNWINDOWED_204,UNWINDOWED_205,UNWINDOWED_206,UNWINDOWED_207,UNWINDOWED_208,UNWINDOWED_209,UNWINDOWED_210,UNWINDOWED_211,UNWINDOWED_212,UNWINDOWED_213,UNWINDOWED_214,UNWINDOWED_215,UNWINDOWED_216,UNWINDOWED_217,UNWINDOWED_218,UNWINDOWED_219,UNWINDOWED_220,UNWINDOWED_221,UNWINDOWED_222,UNWINDOWED_223,UNWINDOWED_224,UNWINDOWED_225,UNWINDOWED_226,UNWINDOWED_227,UNWINDOWED_228,UNWINDOWED_229,UNWINDOWED_230,UNWINDOWED_231,UNWINDOWED_232,UNWINDOWED_233,UNWINDOWED_234,UNWINDOWED_235,UNWINDOWED_236,UNWINDOWED_237,UNWINDOWED_238,UNWINDOWED_239,UNWINDOWED_240,UNWINDOWED_241,UNWINDOWED_242,UNWINDOWED_243,UNWINDOWED_244,UNWINDOWED_245,UNWINDOWED_246,UNWINDOWED_247,UNWINDOWED_248,UNWINDOWED_249,UNWINDOWED_250,UNWINDOWED_251,UNWINDOWED_252,UNWINDOWED_253,UNWINDOWED_254,UNWINDOWED_255,UNWINDOWED_256,UNWINDOWED_257,UNWINDOWED_258,UNWINDOWED_259,UNWINDOWED_260,UNWINDOWED_261,UNWINDOWED_262,UNWINDOWED_263,UNWINDOWED_264,UNWINDOWED_265,UNWINDOWED_266,UNWINDOWED_267,UNWINDOWED_268,UNWINDOWED_269,UNWINDOWED_270,UNWINDOWED_271,UNWINDOWED_272,UNWINDOWED_273,UNWINDOWED_274,UNWINDOWED_275,UNWINDOWED_276,UNWINDOWED_277,UNWINDOWED_278,UNWINDOWED_279,UNWINDOWED_280,UNWINDOWED_281,UNWINDOWED_282,UNWINDOWED_283,UNWINDOWED_284,UNWINDOWED_285,UNWINDOWED_286,UNWINDOWED_287,UNWINDOWED_288,UNWINDOWED_289,UNWINDOWED_290,UNWINDOWED_291,UNWINDOWED_292,UNWINDOWED_293,UNWINDOWED_294,UNWINDOWED_295,UNWINDOWED_296,UNWINDOWED_297,UNWINDOWED_298,UNWINDOWED_299,UNWINDOWED_300,UNWINDOWED_301,UNWINDOWED_302,UNWINDOWED_303,UNWINDOWED_304,UNWINDOWED_305,UNWINDOWED_306,UNWINDOWED_307,UNWINDOWED_308,UNWINDOWED_309,UNWINDOWED_310,UNWINDOWED_311,UNWINDOWED_312,UNWINDOWED_313,UNWINDOWED_314,UNWINDOWED_315,UNWINDOWED_316,UNWINDOWED_317,UNWINDOWED_318,UNWINDOWED_319,UNWINDOWED_320,UNWINDOWED_321,UNWINDOWED_322,UNWINDOWED_323,UNWINDOWED_324,UNWINDOWED_325,UNWINDOWED_326,UNWINDOWED_327,UNWINDOWED_328,UNWINDOWED_329,UNWINDOWED_330,UNWINDOWED_331,UNWINDOWED_332,UNWINDOWED_333,UNWINDOWED_334,UNWINDOWED_335,UNWINDOWED_336,UNWINDOWED_337,UNWINDOWED_338,UNWINDOWED_339,UNWINDOWED_340,UNWINDOWED_341,UNWINDOWED_342,UNWINDOWED_343,UNWINDOWED_344,UNWINDOWED_345,UNWINDOWED_346,UNWINDOWED_347,UNWINDOWED_348,UNWINDOWED_349,UNWINDOWED_350,UNWINDOWED_351,UNWINDOWED_352,UNWINDOWED_353,UNWINDOWED_354,UNWINDOWED_355,UNWINDOWED_356,UNWINDOWED_357,UNWINDOWED_358,UNWINDOWED_359,UNWINDOWED_360,UNWINDOWED_361,UNWINDOWED_362,UNWINDOWED_363,UNWINDOWED_364,UNWINDOWED_365,UNWINDOWED_366,UNWINDOWED_367,UNWINDOWED_368,UNWINDOWED_369,UNWINDOWED_370,UNWINDOWED_371,UNWINDOWED_372,UNWINDOWED_373,UNWINDOWED_374,UNWINDOWED_375,UNWINDOWED_376,UNWINDOWED_377,UNWINDOWED_378,UNWINDOWED_379,UNWINDOWED_380,UNWINDOWED_381,UNWINDOWED_382,UNWINDOWED_383,UNWINDOWED_384,UNWINDOWED_385,UNWINDOWED_386,UNWINDOWED_387,UNWINDOWED_388,UNWINDOWED_389,UNWINDOWED_390,UNWINDOWED_391,UNWINDOWED_392,UNWINDOWED_393,UNWINDOWED_394,UNWINDOWED_395,UNWINDOWED_396,UNWINDOWED_397,UNWINDOWED_398,UNWINDOWED_399,UNWINDOWED_400,UNWINDOWED_401,UNWINDOWED_402,UNWINDOWED_403,UNWINDOWED_404,UNWINDOWED_405,UNWINDOWED_406,UNWINDOWED_407,UNWINDOWED_408,UNWINDOWED_409,UNWINDOWED_410,UNWINDOWED_411,UNWINDOWED_412,UNWINDOWED_413,UNWINDOWED_414,UNWINDOWED_415,UNWINDOWED_416,UNWINDOWED_417,UNWINDOWED_418,UNWINDOWED_419,UNWINDOWED_420,UNWINDOWED_421,UNWINDOWED_422,UNWINDOWED_423,UNWINDOWED_424,UNWINDOWED_425,UNWINDOWED_426,UNWINDOWED_427,UNWINDOWED_428,UNWINDOWED_429,UNWINDOWED_430,UNWINDOWED_431,UNWINDOWED_432,UNWINDOWED_433,UNWINDOWED_434,UNWINDOWED_435,UNWINDOWED_436,UNWINDOWED_437,UNWINDOWED_438,UNWINDOWED_439,UNWINDOWED_440,UNWINDOWED_441,UNWINDOWED_442,UNWINDOWED_443,UNWINDOWED_444,UNWINDOWED_445,UNWINDOWED_446,UNWINDOWED_447,UNWINDOWED_448,UNWINDOWED_449,UNWINDOWED_450,UNWINDOWED_451,UNWINDOWED_452,UNWINDOWED_453,UNWINDOWED_454,UNWINDOWED_455,UNWINDOWED_456,UNWINDOWED_457,UNWINDOWED_458,UNWINDOWED_459,UNWINDOWED_460,UNWINDOWED_461,UNWINDOWED_462,UNWINDOWED_463,UNWINDOWED_464,UNWINDOWED_465,UNWINDOWED_466,UNWINDOWED_467,UNWINDOWED_468,UNWINDOWED_469,UNWINDOWED_470,UNWINDOWED_471,UNWINDOWED_472,UNWINDOWED_473,UNWINDOWED_474,UNWINDOWED_475,UNWINDOWED_476,UNWINDOWED_477,UNWINDOWED_478,UNWINDOWED_479,UNWINDOWED_480,UNWINDOWED_481,UNWINDOWED_482,UNWINDOWED_483,UNWINDOWED_484,UNWINDOWED_485,UNWINDOWED_486,UNWINDOWED_487,UNWINDOWED_488,UNWINDOWED_489,UNWINDOWED_490,UNWINDOWED_491,UNWINDOWED_492,UNWINDOWED_493,UNWINDOWED_494,UNWINDOWED_495,UNWINDOWED_496,UNWINDOWED_497,UNWINDOWED_498,UNWINDOWED_499,UNWINDOWED_500,UNWINDOWED_501,UNWINDOWED_502,UNWINDOWED_503,UNWINDOWED_504,UNWINDOWED_505,UNWINDOWED_506,UNWINDOWED_507,UNWINDOWED_508,UNWINDOWED_509,UNWINDOWED_510,UNWINDOWED_511,UNWINDOWED_512,UNWINDOWED_513,UNWINDOWED_514,UNWINDOWED_515,UNWINDOWED_516,UNWINDOWED_517,UNWINDOWED_518,UNWINDOWED_519,UNWINDOWED_520,UNWINDOWED_521,UNWINDOWED_522,UNWINDOWED_523,UNWINDOWED_524,UNWINDOWED_525,UNWINDOWED_526,UNWINDOWED_527,UNWINDOWED_528,UNWINDOWED_529,UNWINDOWED_530,UNWINDOWED_531,UNWINDOWED_532,UNWINDOWED_533,UNWINDOWED_534,UNWINDOWED_535,UNWINDOWED_536,UNWINDOWED_537,UNWINDOWED_538,UNWINDOWED_539,UNWINDOWED_540,UNWINDOWED_541,UNWINDOWED_542,UNWINDOWED_543,UNWINDOWED_544,UNWINDOWED_545,UNWINDOWED_546,UNWINDOWED_547,UNWINDOWED_548,UNWINDOWED_549,UNWINDOWED_550,UNWINDOWED_551,UNWINDOWED_552,UNWINDOWED_553,UNWINDOWED_554,UNWINDOWED_555,UNWINDOWED_556,UNWINDOWED_557,UNWINDOWED_558,UNWINDOWED_559,UNWINDOWED_560,UNWINDOWED_561,UNWINDOWED_562,UNWINDOWED_563,UNWINDOWED_564,UNWINDOWED_565,UNWINDOWED_566,UNWINDOWED_567,UNWINDOWED_568,UNWINDOWED_569,UNWINDOWED_570,UNWINDOWED_571,UNWINDOWED_572,UNWINDOWED_573,UNWINDOWED_574,UNWINDOWED_575,UNWINDOWED_576,UNWINDOWED_577,UNWINDOWED_578,UNWINDOWED_579,UNWINDOWED_580,UNWINDOWED_581,UNWINDOWED_582,UNWINDOWED_583,UNWINDOWED_584,UNWINDOWED_585,UNWINDOWED_586,UNWINDOWED_587,UNWINDOWED_588,UNWINDOWED_589,UNWINDOWED_590,UNWINDOWED_591,UNWINDOWED_592,UNWINDOWED_593,UNWINDOWED_594,UNWINDOWED_595,UNWINDOWED_596,UNWINDOWED_597,UNWINDOWED_598,UNWINDOWED_599,UNWINDOWED_600,UNWINDOWED_601,UNWINDOWED_602,UNWINDOWED_603,UNWINDOWED_604,UNWINDOWED_605,UNWINDOWED_606,UNWINDOWED_607,UNWINDOWED_608,UNWINDOWED_609,UNWINDOWED_610,UNWINDOWED_611,UNWINDOWED_612,UNWINDOWED_613,UNWINDOWED_614,UNWINDOWED_615,UNWINDOWED_616,UNWINDOWED_617,UNWINDOWED_618,UNWINDOWED_619,UNWINDOWED_620,UNWINDOWED_621,UNWINDOWED_622,UNWINDOWED_623,UNWINDOWED_624,UNWINDOWED_625,UNWINDOWED_626,UNWINDOWED_627,UNWINDOWED_628,UNWINDOWED_629,UNWINDOWED_630,UNWINDOWED_631,UNWINDOWED_632,UNWINDOWED_633,UNWINDOWED_634,UNWINDOWED_635,UNWINDOWED_636,UNWINDOWED_637,UNWINDOWED_638,UNWINDOWED_639,UNWINDOWED_640,UNWINDOWED_641,UNWINDOWED_642,UNWINDOWED_643,UNWINDOWED_644,UNWINDOWED_645,UNWINDOWED_646,UNWINDOWED_647,UNWINDOWED_648,UNWINDOWED_649,UNWINDOWED_650,UNWINDOWED_651,UNWINDOWED_652,UNWINDOWED_653,UNWINDOWED_654,UNWINDOWED_655,UNWINDOWED_656,UNWINDOWED_657,UNWINDOWED_658,UNWINDOWED_659,UNWINDOWED_660,UNWINDOWED_661,UNWINDOWED_662,UNWINDOWED_663,UNWINDOWED_664,UNWINDOWED_665,UNWINDOWED_666,UNWINDOWED_667,UNWINDOWED_668,UNWINDOWED_669,UNWINDOWED_670,UNWINDOWED_671,UNWINDOWED_672,UNWINDOWED_673,UNWINDOWED_674,UNWINDOWED_675,UNWINDOWED_676,UNWINDOWED_677,UNWINDOWED_678,UNWINDOWED_679,UNWINDOWED_680,UNWINDOWED_681,UNWINDOWED_682,UNWINDOWED_683,UNWINDOWED_684,UNWINDOWED_685,UNWINDOWED_686,UNWINDOWED_687,UNWINDOWED_688,UNWINDOWED_689,UNWINDOWED_690,UNWINDOWED_691,UNWINDOWED_692,UNWINDOWED_693,UNWINDOWED_694,UNWINDOWED_695,UNWINDOWED_696,UNWINDOWED_697,UNWINDOWED_698,UNWINDOWED_699,UNWINDOWED_700,UNWINDOWED_701,UNWINDOWED_702,UNWINDOWED_703,UNWINDOWED_704,UNWINDOWED_705,UNWINDOWED_706,UNWINDOWED_707,UNWINDOWED_708,UNWINDOWED_709,UNWINDOWED_710,UNWINDOWED_711,UNWINDOWED_712,UNWINDOWED_713,UNWINDOWED_714,UNWINDOWED_715,UNWINDOWED_716,UNWINDOWED_717,UNWINDOWED_718,UNWINDOWED_719,UNWINDOWED_720,UNWINDOWED_721,UNWINDOWED_722,UNWINDOWED_723,UNWINDOWED_724,UNWINDOWED_725,UNWINDOWED_726,UNWINDOWED_727,UNWINDOWED_728,UNWINDOWED_729,UNWINDOWED_730,UNWINDOWED_731,UNWINDOWED_732,UNWINDOWED_733,UNWINDOWED_734,UNWINDOWED_735,UNWINDOWED_736,UNWINDOWED_737,UNWINDOWED_738,UNWINDOWED_739,UNWINDOWED_740,UNWINDOWED_741,UNWINDOWED_742,UNWINDOWED_743,UNWINDOWED_744,UNWINDOWED_745,UNWINDOWED_746,UNWINDOWED_747,UNWINDOWED_748,UNWINDOWED_749,UNWINDOWED_750,UNWINDOWED_751,UNWINDOWED_752,UNWINDOWED_753,UNWINDOWED_754,UNWINDOWED_755,UNWINDOWED_756,UNWINDOWED_757,UNWINDOWED_758,UNWINDOWED_759,UNWINDOWED_760,UNWINDOWED_761,UNWINDOWED_762,UNWINDOWED_763,UNWINDOWED_764,UNWINDOWED_765,UNWINDOWED_766,UNWINDOWED_767,UNWINDOWED_768,UNWINDOWED_769,UNWINDOWED_770,UNWINDOWED_771,UNWINDOWED_772,UNWINDOWED_773,UNWINDOWED_774,UNWINDOWED_775,UNWINDOWED_776,UNWINDOWED_777,UNWINDOWED_778,UNWINDOWED_779,UNWINDOWED_780,UNWINDOWED_781,UNWINDOWED_782,UNWINDOWED_783,UNWINDOWED_784,UNWINDOWED_785,UNWINDOWED_786,UNWINDOWED_787,UNWINDOWED_788,UNWINDOWED_789,UNWINDOWED_790,UNWINDOWED_791,UNWINDOWED_792,UNWINDOWED_793,UNWINDOWED_794,UNWINDOWED_795,UNWINDOWED_796,UNWINDOWED_797,UNWINDOWED_798,UNWINDOWED_799,UNWINDOWED_800,UNWINDOWED_801,UNWINDOWED_802,UNWINDOWED_803,UNWINDOWED_804,UNWINDOWED_805,UNWINDOWED_806,UNWINDOWED_807,UNWINDOWED_808,UNWINDOWED_809,UNWINDOWED_810,UNWINDOWED_811,UNWINDOWED_812,UNWINDOWED_813,UNWINDOWED_814,UNWINDOWED_815,UNWINDOWED_816,UNWINDOWED_817,UNWINDOWED_818,UNWINDOWED_819,UNWINDOWED_820,UNWINDOWED_821,UNWINDOWED_822,UNWINDOWED_823,UNWINDOWED_824,UNWINDOWED_825,UNWINDOWED_826,UNWINDOWED_827,UNWINDOWED_828,UNWINDOWED_829,UNWINDOWED_830,UNWINDOWED_831,UNWINDOWED_832,UNWINDOWED_833,UNWINDOWED_834,UNWINDOWED_835,UNWINDOWED_836,UNWINDOWED_837,UNWINDOWED_838,UNWINDOWED_839,UNWINDOWED_840,UNWINDOWED_841,UNWINDOWED_842,UNWINDOWED_843,UNWINDOWED_844,UNWINDOWED_845,UNWINDOWED_846,UNWINDOWED_847,UNWINDOWED_848,UNWINDOWED_849,UNWINDOWED_850,UNWINDOWED_851,UNWINDOWED_852,UNWINDOWED_853,UNWINDOWED_854,UNWINDOWED_855,UNWINDOWED_856,UNWINDOWED_857,UNWINDOWED_858,UNWINDOWED_859,UNWINDOWED_860,UNWINDOWED_861,UNWINDOWED_862,UNWINDOWED_863,UNWINDOWED_864,UNWINDOWED_865,UNWINDOWED_866,UNWINDOWED_867,UNWINDOWED_868,UNWINDOWED_869,UNWINDOWED_870,UNWINDOWED_871,UNWINDOWED_872,UNWINDOWED_873,UNWINDOWED_874,UNWINDOWED_875,UNWINDOWED_876,UNWINDOWED_877,UNWINDOWED_878,UNWINDOWED_879,UNWINDOWED_880,UNWINDOWED_881,UNWINDOWED_882,UNWINDOWED_883,UNWINDOWED_884,UNWINDOWED_885,UNWINDOWED_886,UNWINDOWED_887,UNWINDOWED_888,UNWINDOWED_889,UNWINDOWED_890,UNWINDOWED_891,UNWINDOWED_892,UNWINDOWED_893,UNWINDOWED_894,UNWINDOWED_895,UNWINDOWED_896,UNWINDOWED_897,UNWINDOWED_898,UNWINDOWED_899,UNWINDOWED_900,UNWINDOWED_901,UNWINDOWED_902,UNWINDOWED_903,UNWINDOWED_904,UNWINDOWED_905,UNWINDOWED_906,UNWINDOWED_907,UNWINDOWED_908,UNWINDOWED_909,UNWINDOWED_910,UNWINDOWED_911,UNWINDOWED_912,UNWINDOWED_913,UNWINDOWED_914,UNWINDOWED_915,UNWINDOWED_916,UNWINDOWED_917,UNWINDOWED_918,UNWINDOWED_919,UNWINDOWED_920,UNWINDOWED_921,UNWINDOWED_922,UNWINDOWED_923,UNWINDOWED_924,UNWINDOWED_925,UNWINDOWED_926,UNWINDOWED_927,UNWINDOWED_928,UNWINDOWED_929,UNWINDOWED_930,UNWINDOWED_931,UNWINDOWED_932,UNWINDOWED_933,UNWINDOWED_934,UNWINDOWED_935,UNWINDOWED_936,UNWINDOWED_937,UNWINDOWED_938,UNWINDOWED_939,UNWINDOWED_940,UNWINDOWED_941,UNWINDOWED_942,UNWINDOWED_943,UNWINDOWED_944,UNWINDOWED_945,UNWINDOWED_946,UNWINDOWED_947,UNWINDOWED_948,UNWINDOWED_949,UNWINDOWED_950,UNWINDOWED_951,UNWINDOWED_952,UNWINDOWED_953,UNWINDOWED_954,UNWINDOWED_955,UNWINDOWED_956,UNWINDOWED_957,UNWINDOWED_958,UNWINDOWED_959,UNWINDOWED_960,UNWINDOWED_961,UNWINDOWED_962,UNWINDOWED_963,UNWINDOWED_964,UNWINDOWED_965,UNWINDOWED_966,UNWINDOWED_967,UNWINDOWED_968,UNWINDOWED_969,UNWINDOWED_970,UNWINDOWED_971,UNWINDOWED_972,UNWINDOWED_973,UNWINDOWED_974,UNWINDOWED_975,UNWINDOWED_976,UNWINDOWED_977,UNWINDOWED_978,UNWINDOWED_979,UNWINDOWED_980,UNWINDOWED_981,UNWINDOWED_982,UNWINDOWED_983,UNWINDOWED_984,UNWINDOWED_985,UNWINDOWED_986,UNWINDOWED_987,UNWINDOWED_988,UNWINDOWED_989,UNWINDOWED_990,UNWINDOWED_991,UNWINDOWED_992,UNWINDOWED_993,UNWINDOWED_994,UNWINDOWED_995,UNWINDOWED_996,UNWINDOWED_997,UNWINDOWED_998,UNWINDOWED_999,UNWINDOWED_1000,UNWINDOWED_1001,UNWINDOWED_1002,UNWINDOWED_1003,UNWINDOWED_1004,UNWINDOWED_1005,UNWINDOWED_1006,UNWINDOWED_1007,UNWINDOWED_1008,UNWINDOWED_1009,UNWINDOWED_1010,UNWINDOWED_1011,UNWINDOWED_1012,UNWINDOWED_1013,UNWINDOWED_1014,UNWINDOWED_1015,UNWINDOWED_1016,UNWINDOWED_1017,UNWINDOWED_1018,UNWINDOWED_1019,UNWINDOWED_1020,UNWINDOWED_1021,UNWINDOWED_1022,UNWINDOWED_1023: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_DEC_MASK : STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL UNWINDOWED_MASK, REORDERED_MASK, STATE_UPDATE_MASK : STD_LOGIC_VECTOR(1023 DOWNTO 0);
SIGNAL SELECTED_OUTPUT: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_FIRST_CU_DONE : STD_LOGIC;

BEGIN

STATE_REG_0 : n_bit_register_clear_1
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_0 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(0) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_0);
STATE_REG_1 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1);
STATE_REG_2 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_2 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(2) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_2);
STATE_REG_3 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_3 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(3) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_3);
STATE_REG_4 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_4 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(4) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_4);
STATE_REG_5 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_5 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(5) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_5);
STATE_REG_6 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_6 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(6) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_6);
STATE_REG_7 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_7 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(7) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_7);
STATE_REG_8 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_8 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(8) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_8);
STATE_REG_9 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_9 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(9) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_9);
STATE_REG_10 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_10 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(10) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_10);
STATE_REG_11 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_11 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(11) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_11);
STATE_REG_12 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_12 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(12) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_12);
STATE_REG_13 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_13 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(13) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_13);
STATE_REG_14 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_14 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(14) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_14);
STATE_REG_15 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_15 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(15) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_15);
STATE_REG_16 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_16 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(16) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_16);
STATE_REG_17 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_17 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(17) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_17);
STATE_REG_18 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_18 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(18) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_18);
STATE_REG_19 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_19 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(19) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_19);
STATE_REG_20 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_20 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(20) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_20);
STATE_REG_21 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_21 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(21) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_21);
STATE_REG_22 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_22 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(22) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_22);
STATE_REG_23 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_23 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(23) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_23);
STATE_REG_24 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_24 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(24) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_24);
STATE_REG_25 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_25 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(25) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_25);
STATE_REG_26 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_26 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(26) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_26);
STATE_REG_27 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_27 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(27) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_27);
STATE_REG_28 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_28 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(28) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_28);
STATE_REG_29 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_29 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(29) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_29);
STATE_REG_30 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_30 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(30) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_30);
STATE_REG_31 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_31 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(31) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_31);
STATE_REG_32 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_32 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(32) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_32);
STATE_REG_33 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_33 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(33) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_33);
STATE_REG_34 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_34 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(34) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_34);
STATE_REG_35 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_35 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(35) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_35);
STATE_REG_36 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_36 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(36) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_36);
STATE_REG_37 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_37 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(37) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_37);
STATE_REG_38 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_38 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(38) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_38);
STATE_REG_39 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_39 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(39) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_39);
STATE_REG_40 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_40 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(40) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_40);
STATE_REG_41 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_41 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(41) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_41);
STATE_REG_42 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_42 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(42) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_42);
STATE_REG_43 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_43 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(43) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_43);
STATE_REG_44 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_44 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(44) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_44);
STATE_REG_45 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_45 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(45) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_45);
STATE_REG_46 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_46 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(46) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_46);
STATE_REG_47 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_47 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(47) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_47);
STATE_REG_48 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_48 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(48) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_48);
STATE_REG_49 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_49 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(49) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_49);
STATE_REG_50 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_50 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(50) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_50);
STATE_REG_51 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_51 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(51) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_51);
STATE_REG_52 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_52 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(52) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_52);
STATE_REG_53 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_53 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(53) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_53);
STATE_REG_54 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_54 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(54) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_54);
STATE_REG_55 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_55 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(55) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_55);
STATE_REG_56 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_56 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(56) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_56);
STATE_REG_57 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_57 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(57) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_57);
STATE_REG_58 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_58 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(58) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_58);
STATE_REG_59 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_59 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(59) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_59);
STATE_REG_60 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_60 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(60) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_60);
STATE_REG_61 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_61 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(61) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_61);
STATE_REG_62 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_62 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(62) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_62);
STATE_REG_63 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_63 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(63) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_63);
STATE_REG_64 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_64 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(64) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_64);
STATE_REG_65 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_65 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(65) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_65);
STATE_REG_66 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_66 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(66) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_66);
STATE_REG_67 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_67 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(67) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_67);
STATE_REG_68 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_68 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(68) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_68);
STATE_REG_69 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_69 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(69) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_69);
STATE_REG_70 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_70 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(70) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_70);
STATE_REG_71 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_71 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(71) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_71);
STATE_REG_72 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_72 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(72) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_72);
STATE_REG_73 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_73 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(73) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_73);
STATE_REG_74 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_74 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(74) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_74);
STATE_REG_75 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_75 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(75) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_75);
STATE_REG_76 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_76 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(76) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_76);
STATE_REG_77 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_77 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(77) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_77);
STATE_REG_78 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_78 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(78) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_78);
STATE_REG_79 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_79 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(79) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_79);
STATE_REG_80 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_80 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(80) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_80);
STATE_REG_81 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_81 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(81) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_81);
STATE_REG_82 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_82 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(82) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_82);
STATE_REG_83 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_83 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(83) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_83);
STATE_REG_84 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_84 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(84) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_84);
STATE_REG_85 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_85 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(85) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_85);
STATE_REG_86 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_86 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(86) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_86);
STATE_REG_87 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_87 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(87) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_87);
STATE_REG_88 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_88 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(88) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_88);
STATE_REG_89 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_89 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(89) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_89);
STATE_REG_90 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_90 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(90) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_90);
STATE_REG_91 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_91 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(91) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_91);
STATE_REG_92 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_92 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(92) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_92);
STATE_REG_93 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_93 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(93) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_93);
STATE_REG_94 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_94 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(94) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_94);
STATE_REG_95 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_95 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(95) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_95);
STATE_REG_96 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_96 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(96) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_96);
STATE_REG_97 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_97 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(97) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_97);
STATE_REG_98 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_98 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(98) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_98);
STATE_REG_99 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_99 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(99) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_99);
STATE_REG_100 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_100 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(100) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_100);
STATE_REG_101 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_101 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(101) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_101);
STATE_REG_102 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_102 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(102) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_102);
STATE_REG_103 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_103 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(103) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_103);
STATE_REG_104 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_104 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(104) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_104);
STATE_REG_105 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_105 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(105) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_105);
STATE_REG_106 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_106 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(106) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_106);
STATE_REG_107 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_107 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(107) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_107);
STATE_REG_108 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_108 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(108) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_108);
STATE_REG_109 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_109 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(109) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_109);
STATE_REG_110 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_110 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(110) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_110);
STATE_REG_111 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_111 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(111) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_111);
STATE_REG_112 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_112 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(112) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_112);
STATE_REG_113 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_113 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(113) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_113);
STATE_REG_114 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_114 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(114) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_114);
STATE_REG_115 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_115 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(115) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_115);
STATE_REG_116 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_116 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(116) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_116);
STATE_REG_117 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_117 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(117) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_117);
STATE_REG_118 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_118 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(118) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_118);
STATE_REG_119 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_119 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(119) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_119);
STATE_REG_120 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_120 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(120) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_120);
STATE_REG_121 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_121 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(121) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_121);
STATE_REG_122 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_122 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(122) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_122);
STATE_REG_123 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_123 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(123) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_123);
STATE_REG_124 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_124 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(124) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_124);
STATE_REG_125 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_125 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(125) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_125);
STATE_REG_126 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_126 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(126) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_126);
STATE_REG_127 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_127 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(127) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_127);
STATE_REG_128 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_128 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(128) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_128);
STATE_REG_129 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_129 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(129) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_129);
STATE_REG_130 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_130 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(130) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_130);
STATE_REG_131 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_131 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(131) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_131);
STATE_REG_132 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_132 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(132) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_132);
STATE_REG_133 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_133 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(133) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_133);
STATE_REG_134 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_134 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(134) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_134);
STATE_REG_135 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_135 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(135) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_135);
STATE_REG_136 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_136 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(136) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_136);
STATE_REG_137 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_137 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(137) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_137);
STATE_REG_138 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_138 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(138) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_138);
STATE_REG_139 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_139 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(139) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_139);
STATE_REG_140 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_140 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(140) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_140);
STATE_REG_141 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_141 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(141) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_141);
STATE_REG_142 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_142 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(142) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_142);
STATE_REG_143 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_143 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(143) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_143);
STATE_REG_144 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_144 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(144) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_144);
STATE_REG_145 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_145 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(145) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_145);
STATE_REG_146 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_146 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(146) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_146);
STATE_REG_147 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_147 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(147) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_147);
STATE_REG_148 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_148 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(148) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_148);
STATE_REG_149 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_149 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(149) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_149);
STATE_REG_150 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_150 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(150) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_150);
STATE_REG_151 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_151 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(151) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_151);
STATE_REG_152 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_152 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(152) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_152);
STATE_REG_153 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_153 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(153) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_153);
STATE_REG_154 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_154 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(154) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_154);
STATE_REG_155 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_155 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(155) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_155);
STATE_REG_156 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_156 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(156) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_156);
STATE_REG_157 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_157 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(157) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_157);
STATE_REG_158 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_158 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(158) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_158);
STATE_REG_159 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_159 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(159) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_159);
STATE_REG_160 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_160 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(160) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_160);
STATE_REG_161 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_161 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(161) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_161);
STATE_REG_162 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_162 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(162) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_162);
STATE_REG_163 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_163 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(163) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_163);
STATE_REG_164 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_164 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(164) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_164);
STATE_REG_165 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_165 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(165) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_165);
STATE_REG_166 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_166 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(166) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_166);
STATE_REG_167 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_167 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(167) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_167);
STATE_REG_168 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_168 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(168) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_168);
STATE_REG_169 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_169 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(169) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_169);
STATE_REG_170 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_170 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(170) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_170);
STATE_REG_171 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_171 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(171) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_171);
STATE_REG_172 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_172 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(172) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_172);
STATE_REG_173 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_173 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(173) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_173);
STATE_REG_174 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_174 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(174) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_174);
STATE_REG_175 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_175 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(175) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_175);
STATE_REG_176 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_176 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(176) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_176);
STATE_REG_177 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_177 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(177) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_177);
STATE_REG_178 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_178 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(178) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_178);
STATE_REG_179 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_179 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(179) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_179);
STATE_REG_180 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_180 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(180) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_180);
STATE_REG_181 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_181 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(181) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_181);
STATE_REG_182 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_182 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(182) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_182);
STATE_REG_183 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_183 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(183) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_183);
STATE_REG_184 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_184 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(184) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_184);
STATE_REG_185 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_185 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(185) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_185);
STATE_REG_186 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_186 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(186) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_186);
STATE_REG_187 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_187 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(187) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_187);
STATE_REG_188 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_188 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(188) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_188);
STATE_REG_189 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_189 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(189) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_189);
STATE_REG_190 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_190 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(190) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_190);
STATE_REG_191 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_191 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(191) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_191);
STATE_REG_192 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_192 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(192) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_192);
STATE_REG_193 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_193 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(193) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_193);
STATE_REG_194 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_194 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(194) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_194);
STATE_REG_195 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_195 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(195) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_195);
STATE_REG_196 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_196 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(196) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_196);
STATE_REG_197 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_197 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(197) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_197);
STATE_REG_198 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_198 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(198) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_198);
STATE_REG_199 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_199 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(199) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_199);
STATE_REG_200 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_200 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(200) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_200);
STATE_REG_201 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_201 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(201) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_201);
STATE_REG_202 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_202 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(202) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_202);
STATE_REG_203 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_203 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(203) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_203);
STATE_REG_204 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_204 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(204) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_204);
STATE_REG_205 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_205 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(205) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_205);
STATE_REG_206 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_206 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(206) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_206);
STATE_REG_207 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_207 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(207) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_207);
STATE_REG_208 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_208 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(208) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_208);
STATE_REG_209 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_209 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(209) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_209);
STATE_REG_210 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_210 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(210) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_210);
STATE_REG_211 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_211 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(211) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_211);
STATE_REG_212 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_212 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(212) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_212);
STATE_REG_213 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_213 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(213) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_213);
STATE_REG_214 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_214 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(214) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_214);
STATE_REG_215 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_215 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(215) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_215);
STATE_REG_216 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_216 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(216) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_216);
STATE_REG_217 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_217 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(217) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_217);
STATE_REG_218 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_218 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(218) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_218);
STATE_REG_219 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_219 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(219) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_219);
STATE_REG_220 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_220 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(220) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_220);
STATE_REG_221 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_221 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(221) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_221);
STATE_REG_222 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_222 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(222) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_222);
STATE_REG_223 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_223 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(223) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_223);
STATE_REG_224 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_224 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(224) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_224);
STATE_REG_225 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_225 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(225) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_225);
STATE_REG_226 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_226 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(226) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_226);
STATE_REG_227 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_227 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(227) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_227);
STATE_REG_228 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_228 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(228) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_228);
STATE_REG_229 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_229 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(229) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_229);
STATE_REG_230 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_230 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(230) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_230);
STATE_REG_231 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_231 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(231) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_231);
STATE_REG_232 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_232 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(232) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_232);
STATE_REG_233 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_233 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(233) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_233);
STATE_REG_234 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_234 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(234) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_234);
STATE_REG_235 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_235 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(235) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_235);
STATE_REG_236 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_236 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(236) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_236);
STATE_REG_237 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_237 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(237) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_237);
STATE_REG_238 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_238 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(238) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_238);
STATE_REG_239 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_239 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(239) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_239);
STATE_REG_240 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_240 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(240) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_240);
STATE_REG_241 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_241 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(241) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_241);
STATE_REG_242 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_242 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(242) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_242);
STATE_REG_243 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_243 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(243) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_243);
STATE_REG_244 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_244 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(244) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_244);
STATE_REG_245 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_245 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(245) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_245);
STATE_REG_246 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_246 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(246) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_246);
STATE_REG_247 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_247 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(247) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_247);
STATE_REG_248 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_248 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(248) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_248);
STATE_REG_249 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_249 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(249) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_249);
STATE_REG_250 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_250 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(250) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_250);
STATE_REG_251 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_251 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(251) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_251);
STATE_REG_252 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_252 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(252) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_252);
STATE_REG_253 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_253 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(253) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_253);
STATE_REG_254 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_254 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(254) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_254);
STATE_REG_255 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_255 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(255) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_255);
STATE_REG_256 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_256 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(256) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_256);
STATE_REG_257 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_257 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(257) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_257);
STATE_REG_258 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_258 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(258) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_258);
STATE_REG_259 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_259 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(259) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_259);
STATE_REG_260 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_260 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(260) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_260);
STATE_REG_261 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_261 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(261) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_261);
STATE_REG_262 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_262 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(262) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_262);
STATE_REG_263 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_263 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(263) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_263);
STATE_REG_264 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_264 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(264) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_264);
STATE_REG_265 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_265 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(265) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_265);
STATE_REG_266 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_266 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(266) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_266);
STATE_REG_267 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_267 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(267) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_267);
STATE_REG_268 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_268 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(268) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_268);
STATE_REG_269 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_269 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(269) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_269);
STATE_REG_270 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_270 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(270) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_270);
STATE_REG_271 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_271 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(271) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_271);
STATE_REG_272 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_272 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(272) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_272);
STATE_REG_273 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_273 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(273) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_273);
STATE_REG_274 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_274 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(274) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_274);
STATE_REG_275 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_275 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(275) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_275);
STATE_REG_276 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_276 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(276) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_276);
STATE_REG_277 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_277 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(277) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_277);
STATE_REG_278 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_278 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(278) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_278);
STATE_REG_279 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_279 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(279) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_279);
STATE_REG_280 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_280 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(280) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_280);
STATE_REG_281 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_281 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(281) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_281);
STATE_REG_282 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_282 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(282) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_282);
STATE_REG_283 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_283 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(283) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_283);
STATE_REG_284 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_284 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(284) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_284);
STATE_REG_285 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_285 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(285) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_285);
STATE_REG_286 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_286 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(286) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_286);
STATE_REG_287 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_287 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(287) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_287);
STATE_REG_288 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_288 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(288) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_288);
STATE_REG_289 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_289 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(289) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_289);
STATE_REG_290 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_290 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(290) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_290);
STATE_REG_291 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_291 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(291) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_291);
STATE_REG_292 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_292 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(292) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_292);
STATE_REG_293 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_293 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(293) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_293);
STATE_REG_294 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_294 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(294) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_294);
STATE_REG_295 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_295 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(295) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_295);
STATE_REG_296 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_296 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(296) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_296);
STATE_REG_297 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_297 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(297) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_297);
STATE_REG_298 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_298 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(298) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_298);
STATE_REG_299 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_299 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(299) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_299);
STATE_REG_300 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_300 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(300) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_300);
STATE_REG_301 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_301 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(301) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_301);
STATE_REG_302 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_302 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(302) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_302);
STATE_REG_303 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_303 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(303) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_303);
STATE_REG_304 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_304 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(304) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_304);
STATE_REG_305 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_305 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(305) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_305);
STATE_REG_306 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_306 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(306) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_306);
STATE_REG_307 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_307 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(307) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_307);
STATE_REG_308 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_308 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(308) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_308);
STATE_REG_309 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_309 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(309) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_309);
STATE_REG_310 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_310 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(310) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_310);
STATE_REG_311 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_311 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(311) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_311);
STATE_REG_312 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_312 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(312) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_312);
STATE_REG_313 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_313 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(313) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_313);
STATE_REG_314 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_314 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(314) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_314);
STATE_REG_315 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_315 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(315) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_315);
STATE_REG_316 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_316 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(316) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_316);
STATE_REG_317 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_317 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(317) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_317);
STATE_REG_318 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_318 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(318) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_318);
STATE_REG_319 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_319 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(319) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_319);
STATE_REG_320 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_320 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(320) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_320);
STATE_REG_321 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_321 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(321) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_321);
STATE_REG_322 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_322 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(322) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_322);
STATE_REG_323 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_323 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(323) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_323);
STATE_REG_324 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_324 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(324) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_324);
STATE_REG_325 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_325 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(325) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_325);
STATE_REG_326 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_326 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(326) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_326);
STATE_REG_327 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_327 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(327) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_327);
STATE_REG_328 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_328 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(328) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_328);
STATE_REG_329 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_329 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(329) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_329);
STATE_REG_330 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_330 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(330) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_330);
STATE_REG_331 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_331 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(331) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_331);
STATE_REG_332 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_332 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(332) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_332);
STATE_REG_333 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_333 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(333) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_333);
STATE_REG_334 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_334 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(334) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_334);
STATE_REG_335 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_335 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(335) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_335);
STATE_REG_336 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_336 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(336) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_336);
STATE_REG_337 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_337 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(337) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_337);
STATE_REG_338 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_338 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(338) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_338);
STATE_REG_339 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_339 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(339) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_339);
STATE_REG_340 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_340 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(340) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_340);
STATE_REG_341 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_341 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(341) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_341);
STATE_REG_342 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_342 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(342) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_342);
STATE_REG_343 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_343 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(343) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_343);
STATE_REG_344 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_344 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(344) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_344);
STATE_REG_345 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_345 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(345) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_345);
STATE_REG_346 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_346 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(346) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_346);
STATE_REG_347 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_347 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(347) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_347);
STATE_REG_348 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_348 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(348) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_348);
STATE_REG_349 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_349 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(349) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_349);
STATE_REG_350 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_350 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(350) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_350);
STATE_REG_351 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_351 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(351) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_351);
STATE_REG_352 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_352 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(352) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_352);
STATE_REG_353 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_353 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(353) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_353);
STATE_REG_354 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_354 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(354) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_354);
STATE_REG_355 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_355 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(355) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_355);
STATE_REG_356 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_356 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(356) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_356);
STATE_REG_357 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_357 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(357) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_357);
STATE_REG_358 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_358 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(358) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_358);
STATE_REG_359 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_359 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(359) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_359);
STATE_REG_360 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_360 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(360) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_360);
STATE_REG_361 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_361 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(361) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_361);
STATE_REG_362 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_362 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(362) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_362);
STATE_REG_363 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_363 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(363) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_363);
STATE_REG_364 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_364 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(364) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_364);
STATE_REG_365 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_365 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(365) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_365);
STATE_REG_366 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_366 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(366) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_366);
STATE_REG_367 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_367 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(367) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_367);
STATE_REG_368 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_368 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(368) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_368);
STATE_REG_369 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_369 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(369) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_369);
STATE_REG_370 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_370 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(370) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_370);
STATE_REG_371 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_371 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(371) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_371);
STATE_REG_372 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_372 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(372) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_372);
STATE_REG_373 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_373 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(373) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_373);
STATE_REG_374 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_374 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(374) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_374);
STATE_REG_375 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_375 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(375) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_375);
STATE_REG_376 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_376 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(376) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_376);
STATE_REG_377 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_377 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(377) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_377);
STATE_REG_378 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_378 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(378) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_378);
STATE_REG_379 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_379 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(379) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_379);
STATE_REG_380 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_380 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(380) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_380);
STATE_REG_381 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_381 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(381) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_381);
STATE_REG_382 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_382 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(382) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_382);
STATE_REG_383 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_383 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(383) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_383);
STATE_REG_384 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_384 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(384) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_384);
STATE_REG_385 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_385 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(385) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_385);
STATE_REG_386 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_386 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(386) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_386);
STATE_REG_387 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_387 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(387) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_387);
STATE_REG_388 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_388 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(388) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_388);
STATE_REG_389 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_389 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(389) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_389);
STATE_REG_390 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_390 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(390) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_390);
STATE_REG_391 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_391 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(391) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_391);
STATE_REG_392 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_392 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(392) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_392);
STATE_REG_393 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_393 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(393) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_393);
STATE_REG_394 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_394 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(394) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_394);
STATE_REG_395 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_395 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(395) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_395);
STATE_REG_396 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_396 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(396) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_396);
STATE_REG_397 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_397 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(397) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_397);
STATE_REG_398 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_398 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(398) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_398);
STATE_REG_399 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_399 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(399) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_399);
STATE_REG_400 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_400 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(400) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_400);
STATE_REG_401 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_401 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(401) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_401);
STATE_REG_402 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_402 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(402) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_402);
STATE_REG_403 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_403 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(403) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_403);
STATE_REG_404 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_404 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(404) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_404);
STATE_REG_405 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_405 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(405) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_405);
STATE_REG_406 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_406 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(406) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_406);
STATE_REG_407 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_407 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(407) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_407);
STATE_REG_408 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_408 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(408) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_408);
STATE_REG_409 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_409 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(409) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_409);
STATE_REG_410 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_410 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(410) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_410);
STATE_REG_411 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_411 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(411) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_411);
STATE_REG_412 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_412 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(412) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_412);
STATE_REG_413 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_413 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(413) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_413);
STATE_REG_414 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_414 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(414) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_414);
STATE_REG_415 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_415 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(415) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_415);
STATE_REG_416 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_416 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(416) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_416);
STATE_REG_417 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_417 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(417) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_417);
STATE_REG_418 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_418 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(418) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_418);
STATE_REG_419 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_419 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(419) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_419);
STATE_REG_420 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_420 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(420) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_420);
STATE_REG_421 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_421 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(421) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_421);
STATE_REG_422 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_422 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(422) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_422);
STATE_REG_423 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_423 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(423) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_423);
STATE_REG_424 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_424 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(424) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_424);
STATE_REG_425 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_425 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(425) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_425);
STATE_REG_426 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_426 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(426) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_426);
STATE_REG_427 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_427 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(427) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_427);
STATE_REG_428 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_428 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(428) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_428);
STATE_REG_429 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_429 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(429) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_429);
STATE_REG_430 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_430 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(430) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_430);
STATE_REG_431 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_431 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(431) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_431);
STATE_REG_432 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_432 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(432) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_432);
STATE_REG_433 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_433 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(433) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_433);
STATE_REG_434 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_434 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(434) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_434);
STATE_REG_435 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_435 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(435) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_435);
STATE_REG_436 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_436 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(436) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_436);
STATE_REG_437 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_437 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(437) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_437);
STATE_REG_438 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_438 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(438) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_438);
STATE_REG_439 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_439 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(439) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_439);
STATE_REG_440 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_440 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(440) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_440);
STATE_REG_441 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_441 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(441) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_441);
STATE_REG_442 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_442 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(442) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_442);
STATE_REG_443 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_443 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(443) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_443);
STATE_REG_444 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_444 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(444) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_444);
STATE_REG_445 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_445 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(445) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_445);
STATE_REG_446 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_446 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(446) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_446);
STATE_REG_447 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_447 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(447) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_447);
STATE_REG_448 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_448 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(448) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_448);
STATE_REG_449 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_449 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(449) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_449);
STATE_REG_450 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_450 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(450) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_450);
STATE_REG_451 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_451 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(451) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_451);
STATE_REG_452 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_452 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(452) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_452);
STATE_REG_453 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_453 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(453) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_453);
STATE_REG_454 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_454 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(454) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_454);
STATE_REG_455 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_455 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(455) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_455);
STATE_REG_456 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_456 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(456) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_456);
STATE_REG_457 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_457 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(457) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_457);
STATE_REG_458 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_458 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(458) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_458);
STATE_REG_459 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_459 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(459) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_459);
STATE_REG_460 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_460 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(460) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_460);
STATE_REG_461 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_461 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(461) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_461);
STATE_REG_462 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_462 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(462) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_462);
STATE_REG_463 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_463 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(463) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_463);
STATE_REG_464 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_464 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(464) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_464);
STATE_REG_465 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_465 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(465) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_465);
STATE_REG_466 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_466 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(466) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_466);
STATE_REG_467 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_467 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(467) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_467);
STATE_REG_468 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_468 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(468) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_468);
STATE_REG_469 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_469 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(469) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_469);
STATE_REG_470 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_470 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(470) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_470);
STATE_REG_471 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_471 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(471) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_471);
STATE_REG_472 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_472 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(472) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_472);
STATE_REG_473 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_473 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(473) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_473);
STATE_REG_474 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_474 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(474) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_474);
STATE_REG_475 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_475 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(475) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_475);
STATE_REG_476 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_476 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(476) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_476);
STATE_REG_477 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_477 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(477) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_477);
STATE_REG_478 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_478 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(478) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_478);
STATE_REG_479 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_479 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(479) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_479);
STATE_REG_480 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_480 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(480) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_480);
STATE_REG_481 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_481 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(481) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_481);
STATE_REG_482 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_482 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(482) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_482);
STATE_REG_483 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_483 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(483) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_483);
STATE_REG_484 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_484 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(484) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_484);
STATE_REG_485 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_485 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(485) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_485);
STATE_REG_486 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_486 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(486) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_486);
STATE_REG_487 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_487 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(487) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_487);
STATE_REG_488 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_488 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(488) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_488);
STATE_REG_489 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_489 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(489) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_489);
STATE_REG_490 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_490 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(490) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_490);
STATE_REG_491 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_491 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(491) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_491);
STATE_REG_492 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_492 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(492) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_492);
STATE_REG_493 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_493 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(493) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_493);
STATE_REG_494 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_494 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(494) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_494);
STATE_REG_495 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_495 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(495) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_495);
STATE_REG_496 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_496 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(496) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_496);
STATE_REG_497 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_497 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(497) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_497);
STATE_REG_498 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_498 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(498) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_498);
STATE_REG_499 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_499 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(499) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_499);
STATE_REG_500 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_500 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(500) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_500);
STATE_REG_501 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_501 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(501) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_501);
STATE_REG_502 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_502 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(502) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_502);
STATE_REG_503 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_503 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(503) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_503);
STATE_REG_504 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_504 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(504) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_504);
STATE_REG_505 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_505 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(505) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_505);
STATE_REG_506 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_506 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(506) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_506);
STATE_REG_507 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_507 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(507) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_507);
STATE_REG_508 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_508 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(508) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_508);
STATE_REG_509 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_509 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(509) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_509);
STATE_REG_510 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_510 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(510) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_510);
STATE_REG_511 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_511 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(511) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_511);
STATE_REG_512 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_512 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(512) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_512);
STATE_REG_513 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_513 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(513) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_513);
STATE_REG_514 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_514 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(514) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_514);
STATE_REG_515 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_515 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(515) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_515);
STATE_REG_516 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_516 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(516) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_516);
STATE_REG_517 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_517 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(517) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_517);
STATE_REG_518 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_518 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(518) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_518);
STATE_REG_519 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_519 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(519) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_519);
STATE_REG_520 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_520 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(520) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_520);
STATE_REG_521 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_521 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(521) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_521);
STATE_REG_522 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_522 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(522) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_522);
STATE_REG_523 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_523 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(523) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_523);
STATE_REG_524 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_524 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(524) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_524);
STATE_REG_525 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_525 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(525) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_525);
STATE_REG_526 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_526 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(526) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_526);
STATE_REG_527 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_527 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(527) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_527);
STATE_REG_528 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_528 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(528) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_528);
STATE_REG_529 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_529 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(529) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_529);
STATE_REG_530 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_530 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(530) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_530);
STATE_REG_531 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_531 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(531) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_531);
STATE_REG_532 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_532 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(532) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_532);
STATE_REG_533 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_533 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(533) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_533);
STATE_REG_534 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_534 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(534) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_534);
STATE_REG_535 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_535 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(535) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_535);
STATE_REG_536 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_536 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(536) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_536);
STATE_REG_537 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_537 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(537) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_537);
STATE_REG_538 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_538 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(538) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_538);
STATE_REG_539 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_539 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(539) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_539);
STATE_REG_540 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_540 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(540) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_540);
STATE_REG_541 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_541 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(541) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_541);
STATE_REG_542 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_542 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(542) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_542);
STATE_REG_543 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_543 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(543) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_543);
STATE_REG_544 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_544 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(544) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_544);
STATE_REG_545 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_545 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(545) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_545);
STATE_REG_546 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_546 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(546) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_546);
STATE_REG_547 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_547 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(547) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_547);
STATE_REG_548 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_548 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(548) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_548);
STATE_REG_549 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_549 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(549) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_549);
STATE_REG_550 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_550 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(550) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_550);
STATE_REG_551 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_551 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(551) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_551);
STATE_REG_552 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_552 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(552) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_552);
STATE_REG_553 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_553 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(553) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_553);
STATE_REG_554 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_554 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(554) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_554);
STATE_REG_555 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_555 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(555) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_555);
STATE_REG_556 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_556 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(556) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_556);
STATE_REG_557 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_557 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(557) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_557);
STATE_REG_558 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_558 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(558) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_558);
STATE_REG_559 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_559 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(559) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_559);
STATE_REG_560 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_560 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(560) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_560);
STATE_REG_561 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_561 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(561) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_561);
STATE_REG_562 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_562 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(562) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_562);
STATE_REG_563 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_563 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(563) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_563);
STATE_REG_564 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_564 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(564) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_564);
STATE_REG_565 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_565 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(565) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_565);
STATE_REG_566 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_566 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(566) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_566);
STATE_REG_567 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_567 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(567) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_567);
STATE_REG_568 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_568 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(568) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_568);
STATE_REG_569 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_569 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(569) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_569);
STATE_REG_570 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_570 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(570) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_570);
STATE_REG_571 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_571 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(571) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_571);
STATE_REG_572 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_572 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(572) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_572);
STATE_REG_573 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_573 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(573) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_573);
STATE_REG_574 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_574 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(574) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_574);
STATE_REG_575 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_575 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(575) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_575);
STATE_REG_576 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_576 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(576) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_576);
STATE_REG_577 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_577 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(577) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_577);
STATE_REG_578 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_578 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(578) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_578);
STATE_REG_579 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_579 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(579) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_579);
STATE_REG_580 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_580 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(580) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_580);
STATE_REG_581 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_581 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(581) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_581);
STATE_REG_582 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_582 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(582) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_582);
STATE_REG_583 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_583 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(583) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_583);
STATE_REG_584 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_584 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(584) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_584);
STATE_REG_585 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_585 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(585) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_585);
STATE_REG_586 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_586 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(586) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_586);
STATE_REG_587 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_587 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(587) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_587);
STATE_REG_588 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_588 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(588) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_588);
STATE_REG_589 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_589 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(589) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_589);
STATE_REG_590 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_590 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(590) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_590);
STATE_REG_591 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_591 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(591) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_591);
STATE_REG_592 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_592 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(592) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_592);
STATE_REG_593 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_593 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(593) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_593);
STATE_REG_594 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_594 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(594) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_594);
STATE_REG_595 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_595 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(595) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_595);
STATE_REG_596 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_596 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(596) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_596);
STATE_REG_597 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_597 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(597) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_597);
STATE_REG_598 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_598 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(598) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_598);
STATE_REG_599 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_599 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(599) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_599);
STATE_REG_600 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_600 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(600) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_600);
STATE_REG_601 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_601 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(601) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_601);
STATE_REG_602 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_602 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(602) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_602);
STATE_REG_603 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_603 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(603) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_603);
STATE_REG_604 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_604 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(604) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_604);
STATE_REG_605 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_605 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(605) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_605);
STATE_REG_606 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_606 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(606) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_606);
STATE_REG_607 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_607 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(607) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_607);
STATE_REG_608 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_608 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(608) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_608);
STATE_REG_609 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_609 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(609) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_609);
STATE_REG_610 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_610 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(610) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_610);
STATE_REG_611 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_611 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(611) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_611);
STATE_REG_612 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_612 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(612) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_612);
STATE_REG_613 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_613 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(613) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_613);
STATE_REG_614 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_614 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(614) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_614);
STATE_REG_615 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_615 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(615) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_615);
STATE_REG_616 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_616 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(616) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_616);
STATE_REG_617 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_617 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(617) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_617);
STATE_REG_618 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_618 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(618) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_618);
STATE_REG_619 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_619 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(619) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_619);
STATE_REG_620 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_620 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(620) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_620);
STATE_REG_621 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_621 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(621) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_621);
STATE_REG_622 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_622 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(622) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_622);
STATE_REG_623 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_623 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(623) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_623);
STATE_REG_624 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_624 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(624) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_624);
STATE_REG_625 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_625 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(625) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_625);
STATE_REG_626 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_626 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(626) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_626);
STATE_REG_627 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_627 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(627) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_627);
STATE_REG_628 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_628 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(628) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_628);
STATE_REG_629 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_629 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(629) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_629);
STATE_REG_630 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_630 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(630) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_630);
STATE_REG_631 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_631 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(631) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_631);
STATE_REG_632 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_632 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(632) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_632);
STATE_REG_633 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_633 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(633) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_633);
STATE_REG_634 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_634 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(634) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_634);
STATE_REG_635 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_635 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(635) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_635);
STATE_REG_636 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_636 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(636) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_636);
STATE_REG_637 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_637 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(637) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_637);
STATE_REG_638 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_638 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(638) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_638);
STATE_REG_639 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_639 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(639) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_639);
STATE_REG_640 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_640 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(640) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_640);
STATE_REG_641 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_641 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(641) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_641);
STATE_REG_642 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_642 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(642) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_642);
STATE_REG_643 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_643 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(643) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_643);
STATE_REG_644 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_644 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(644) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_644);
STATE_REG_645 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_645 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(645) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_645);
STATE_REG_646 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_646 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(646) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_646);
STATE_REG_647 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_647 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(647) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_647);
STATE_REG_648 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_648 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(648) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_648);
STATE_REG_649 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_649 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(649) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_649);
STATE_REG_650 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_650 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(650) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_650);
STATE_REG_651 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_651 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(651) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_651);
STATE_REG_652 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_652 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(652) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_652);
STATE_REG_653 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_653 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(653) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_653);
STATE_REG_654 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_654 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(654) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_654);
STATE_REG_655 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_655 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(655) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_655);
STATE_REG_656 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_656 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(656) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_656);
STATE_REG_657 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_657 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(657) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_657);
STATE_REG_658 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_658 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(658) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_658);
STATE_REG_659 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_659 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(659) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_659);
STATE_REG_660 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_660 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(660) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_660);
STATE_REG_661 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_661 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(661) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_661);
STATE_REG_662 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_662 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(662) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_662);
STATE_REG_663 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_663 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(663) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_663);
STATE_REG_664 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_664 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(664) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_664);
STATE_REG_665 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_665 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(665) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_665);
STATE_REG_666 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_666 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(666) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_666);
STATE_REG_667 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_667 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(667) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_667);
STATE_REG_668 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_668 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(668) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_668);
STATE_REG_669 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_669 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(669) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_669);
STATE_REG_670 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_670 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(670) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_670);
STATE_REG_671 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_671 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(671) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_671);
STATE_REG_672 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_672 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(672) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_672);
STATE_REG_673 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_673 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(673) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_673);
STATE_REG_674 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_674 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(674) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_674);
STATE_REG_675 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_675 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(675) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_675);
STATE_REG_676 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_676 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(676) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_676);
STATE_REG_677 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_677 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(677) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_677);
STATE_REG_678 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_678 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(678) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_678);
STATE_REG_679 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_679 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(679) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_679);
STATE_REG_680 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_680 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(680) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_680);
STATE_REG_681 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_681 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(681) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_681);
STATE_REG_682 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_682 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(682) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_682);
STATE_REG_683 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_683 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(683) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_683);
STATE_REG_684 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_684 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(684) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_684);
STATE_REG_685 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_685 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(685) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_685);
STATE_REG_686 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_686 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(686) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_686);
STATE_REG_687 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_687 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(687) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_687);
STATE_REG_688 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_688 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(688) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_688);
STATE_REG_689 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_689 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(689) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_689);
STATE_REG_690 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_690 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(690) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_690);
STATE_REG_691 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_691 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(691) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_691);
STATE_REG_692 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_692 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(692) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_692);
STATE_REG_693 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_693 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(693) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_693);
STATE_REG_694 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_694 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(694) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_694);
STATE_REG_695 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_695 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(695) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_695);
STATE_REG_696 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_696 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(696) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_696);
STATE_REG_697 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_697 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(697) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_697);
STATE_REG_698 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_698 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(698) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_698);
STATE_REG_699 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_699 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(699) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_699);
STATE_REG_700 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_700 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(700) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_700);
STATE_REG_701 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_701 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(701) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_701);
STATE_REG_702 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_702 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(702) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_702);
STATE_REG_703 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_703 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(703) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_703);
STATE_REG_704 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_704 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(704) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_704);
STATE_REG_705 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_705 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(705) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_705);
STATE_REG_706 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_706 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(706) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_706);
STATE_REG_707 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_707 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(707) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_707);
STATE_REG_708 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_708 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(708) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_708);
STATE_REG_709 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_709 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(709) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_709);
STATE_REG_710 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_710 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(710) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_710);
STATE_REG_711 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_711 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(711) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_711);
STATE_REG_712 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_712 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(712) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_712);
STATE_REG_713 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_713 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(713) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_713);
STATE_REG_714 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_714 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(714) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_714);
STATE_REG_715 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_715 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(715) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_715);
STATE_REG_716 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_716 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(716) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_716);
STATE_REG_717 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_717 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(717) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_717);
STATE_REG_718 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_718 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(718) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_718);
STATE_REG_719 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_719 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(719) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_719);
STATE_REG_720 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_720 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(720) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_720);
STATE_REG_721 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_721 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(721) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_721);
STATE_REG_722 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_722 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(722) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_722);
STATE_REG_723 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_723 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(723) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_723);
STATE_REG_724 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_724 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(724) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_724);
STATE_REG_725 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_725 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(725) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_725);
STATE_REG_726 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_726 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(726) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_726);
STATE_REG_727 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_727 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(727) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_727);
STATE_REG_728 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_728 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(728) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_728);
STATE_REG_729 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_729 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(729) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_729);
STATE_REG_730 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_730 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(730) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_730);
STATE_REG_731 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_731 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(731) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_731);
STATE_REG_732 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_732 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(732) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_732);
STATE_REG_733 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_733 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(733) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_733);
STATE_REG_734 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_734 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(734) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_734);
STATE_REG_735 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_735 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(735) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_735);
STATE_REG_736 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_736 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(736) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_736);
STATE_REG_737 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_737 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(737) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_737);
STATE_REG_738 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_738 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(738) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_738);
STATE_REG_739 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_739 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(739) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_739);
STATE_REG_740 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_740 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(740) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_740);
STATE_REG_741 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_741 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(741) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_741);
STATE_REG_742 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_742 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(742) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_742);
STATE_REG_743 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_743 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(743) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_743);
STATE_REG_744 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_744 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(744) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_744);
STATE_REG_745 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_745 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(745) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_745);
STATE_REG_746 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_746 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(746) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_746);
STATE_REG_747 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_747 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(747) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_747);
STATE_REG_748 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_748 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(748) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_748);
STATE_REG_749 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_749 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(749) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_749);
STATE_REG_750 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_750 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(750) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_750);
STATE_REG_751 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_751 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(751) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_751);
STATE_REG_752 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_752 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(752) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_752);
STATE_REG_753 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_753 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(753) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_753);
STATE_REG_754 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_754 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(754) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_754);
STATE_REG_755 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_755 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(755) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_755);
STATE_REG_756 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_756 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(756) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_756);
STATE_REG_757 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_757 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(757) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_757);
STATE_REG_758 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_758 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(758) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_758);
STATE_REG_759 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_759 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(759) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_759);
STATE_REG_760 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_760 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(760) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_760);
STATE_REG_761 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_761 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(761) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_761);
STATE_REG_762 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_762 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(762) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_762);
STATE_REG_763 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_763 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(763) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_763);
STATE_REG_764 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_764 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(764) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_764);
STATE_REG_765 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_765 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(765) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_765);
STATE_REG_766 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_766 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(766) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_766);
STATE_REG_767 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_767 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(767) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_767);
STATE_REG_768 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_768 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(768) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_768);
STATE_REG_769 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_769 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(769) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_769);
STATE_REG_770 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_770 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(770) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_770);
STATE_REG_771 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_771 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(771) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_771);
STATE_REG_772 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_772 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(772) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_772);
STATE_REG_773 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_773 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(773) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_773);
STATE_REG_774 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_774 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(774) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_774);
STATE_REG_775 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_775 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(775) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_775);
STATE_REG_776 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_776 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(776) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_776);
STATE_REG_777 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_777 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(777) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_777);
STATE_REG_778 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_778 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(778) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_778);
STATE_REG_779 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_779 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(779) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_779);
STATE_REG_780 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_780 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(780) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_780);
STATE_REG_781 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_781 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(781) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_781);
STATE_REG_782 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_782 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(782) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_782);
STATE_REG_783 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_783 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(783) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_783);
STATE_REG_784 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_784 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(784) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_784);
STATE_REG_785 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_785 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(785) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_785);
STATE_REG_786 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_786 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(786) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_786);
STATE_REG_787 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_787 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(787) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_787);
STATE_REG_788 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_788 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(788) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_788);
STATE_REG_789 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_789 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(789) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_789);
STATE_REG_790 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_790 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(790) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_790);
STATE_REG_791 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_791 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(791) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_791);
STATE_REG_792 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_792 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(792) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_792);
STATE_REG_793 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_793 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(793) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_793);
STATE_REG_794 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_794 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(794) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_794);
STATE_REG_795 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_795 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(795) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_795);
STATE_REG_796 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_796 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(796) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_796);
STATE_REG_797 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_797 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(797) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_797);
STATE_REG_798 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_798 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(798) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_798);
STATE_REG_799 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_799 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(799) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_799);
STATE_REG_800 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_800 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(800) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_800);
STATE_REG_801 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_801 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(801) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_801);
STATE_REG_802 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_802 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(802) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_802);
STATE_REG_803 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_803 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(803) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_803);
STATE_REG_804 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_804 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(804) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_804);
STATE_REG_805 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_805 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(805) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_805);
STATE_REG_806 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_806 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(806) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_806);
STATE_REG_807 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_807 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(807) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_807);
STATE_REG_808 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_808 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(808) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_808);
STATE_REG_809 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_809 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(809) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_809);
STATE_REG_810 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_810 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(810) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_810);
STATE_REG_811 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_811 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(811) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_811);
STATE_REG_812 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_812 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(812) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_812);
STATE_REG_813 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_813 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(813) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_813);
STATE_REG_814 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_814 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(814) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_814);
STATE_REG_815 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_815 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(815) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_815);
STATE_REG_816 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_816 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(816) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_816);
STATE_REG_817 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_817 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(817) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_817);
STATE_REG_818 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_818 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(818) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_818);
STATE_REG_819 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_819 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(819) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_819);
STATE_REG_820 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_820 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(820) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_820);
STATE_REG_821 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_821 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(821) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_821);
STATE_REG_822 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_822 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(822) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_822);
STATE_REG_823 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_823 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(823) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_823);
STATE_REG_824 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_824 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(824) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_824);
STATE_REG_825 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_825 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(825) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_825);
STATE_REG_826 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_826 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(826) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_826);
STATE_REG_827 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_827 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(827) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_827);
STATE_REG_828 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_828 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(828) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_828);
STATE_REG_829 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_829 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(829) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_829);
STATE_REG_830 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_830 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(830) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_830);
STATE_REG_831 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_831 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(831) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_831);
STATE_REG_832 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_832 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(832) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_832);
STATE_REG_833 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_833 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(833) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_833);
STATE_REG_834 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_834 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(834) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_834);
STATE_REG_835 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_835 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(835) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_835);
STATE_REG_836 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_836 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(836) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_836);
STATE_REG_837 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_837 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(837) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_837);
STATE_REG_838 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_838 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(838) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_838);
STATE_REG_839 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_839 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(839) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_839);
STATE_REG_840 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_840 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(840) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_840);
STATE_REG_841 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_841 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(841) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_841);
STATE_REG_842 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_842 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(842) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_842);
STATE_REG_843 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_843 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(843) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_843);
STATE_REG_844 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_844 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(844) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_844);
STATE_REG_845 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_845 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(845) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_845);
STATE_REG_846 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_846 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(846) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_846);
STATE_REG_847 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_847 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(847) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_847);
STATE_REG_848 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_848 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(848) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_848);
STATE_REG_849 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_849 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(849) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_849);
STATE_REG_850 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_850 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(850) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_850);
STATE_REG_851 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_851 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(851) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_851);
STATE_REG_852 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_852 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(852) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_852);
STATE_REG_853 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_853 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(853) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_853);
STATE_REG_854 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_854 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(854) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_854);
STATE_REG_855 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_855 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(855) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_855);
STATE_REG_856 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_856 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(856) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_856);
STATE_REG_857 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_857 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(857) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_857);
STATE_REG_858 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_858 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(858) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_858);
STATE_REG_859 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_859 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(859) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_859);
STATE_REG_860 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_860 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(860) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_860);
STATE_REG_861 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_861 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(861) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_861);
STATE_REG_862 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_862 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(862) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_862);
STATE_REG_863 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_863 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(863) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_863);
STATE_REG_864 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_864 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(864) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_864);
STATE_REG_865 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_865 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(865) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_865);
STATE_REG_866 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_866 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(866) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_866);
STATE_REG_867 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_867 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(867) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_867);
STATE_REG_868 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_868 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(868) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_868);
STATE_REG_869 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_869 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(869) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_869);
STATE_REG_870 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_870 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(870) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_870);
STATE_REG_871 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_871 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(871) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_871);
STATE_REG_872 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_872 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(872) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_872);
STATE_REG_873 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_873 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(873) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_873);
STATE_REG_874 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_874 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(874) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_874);
STATE_REG_875 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_875 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(875) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_875);
STATE_REG_876 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_876 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(876) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_876);
STATE_REG_877 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_877 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(877) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_877);
STATE_REG_878 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_878 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(878) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_878);
STATE_REG_879 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_879 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(879) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_879);
STATE_REG_880 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_880 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(880) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_880);
STATE_REG_881 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_881 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(881) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_881);
STATE_REG_882 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_882 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(882) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_882);
STATE_REG_883 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_883 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(883) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_883);
STATE_REG_884 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_884 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(884) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_884);
STATE_REG_885 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_885 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(885) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_885);
STATE_REG_886 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_886 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(886) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_886);
STATE_REG_887 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_887 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(887) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_887);
STATE_REG_888 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_888 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(888) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_888);
STATE_REG_889 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_889 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(889) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_889);
STATE_REG_890 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_890 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(890) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_890);
STATE_REG_891 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_891 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(891) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_891);
STATE_REG_892 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_892 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(892) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_892);
STATE_REG_893 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_893 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(893) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_893);
STATE_REG_894 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_894 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(894) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_894);
STATE_REG_895 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_895 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(895) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_895);
STATE_REG_896 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_896 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(896) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_896);
STATE_REG_897 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_897 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(897) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_897);
STATE_REG_898 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_898 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(898) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_898);
STATE_REG_899 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_899 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(899) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_899);
STATE_REG_900 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_900 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(900) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_900);
STATE_REG_901 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_901 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(901) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_901);
STATE_REG_902 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_902 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(902) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_902);
STATE_REG_903 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_903 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(903) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_903);
STATE_REG_904 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_904 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(904) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_904);
STATE_REG_905 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_905 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(905) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_905);
STATE_REG_906 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_906 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(906) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_906);
STATE_REG_907 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_907 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(907) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_907);
STATE_REG_908 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_908 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(908) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_908);
STATE_REG_909 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_909 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(909) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_909);
STATE_REG_910 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_910 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(910) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_910);
STATE_REG_911 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_911 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(911) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_911);
STATE_REG_912 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_912 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(912) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_912);
STATE_REG_913 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_913 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(913) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_913);
STATE_REG_914 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_914 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(914) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_914);
STATE_REG_915 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_915 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(915) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_915);
STATE_REG_916 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_916 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(916) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_916);
STATE_REG_917 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_917 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(917) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_917);
STATE_REG_918 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_918 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(918) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_918);
STATE_REG_919 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_919 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(919) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_919);
STATE_REG_920 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_920 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(920) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_920);
STATE_REG_921 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_921 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(921) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_921);
STATE_REG_922 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_922 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(922) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_922);
STATE_REG_923 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_923 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(923) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_923);
STATE_REG_924 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_924 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(924) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_924);
STATE_REG_925 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_925 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(925) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_925);
STATE_REG_926 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_926 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(926) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_926);
STATE_REG_927 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_927 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(927) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_927);
STATE_REG_928 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_928 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(928) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_928);
STATE_REG_929 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_929 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(929) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_929);
STATE_REG_930 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_930 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(930) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_930);
STATE_REG_931 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_931 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(931) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_931);
STATE_REG_932 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_932 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(932) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_932);
STATE_REG_933 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_933 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(933) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_933);
STATE_REG_934 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_934 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(934) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_934);
STATE_REG_935 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_935 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(935) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_935);
STATE_REG_936 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_936 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(936) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_936);
STATE_REG_937 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_937 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(937) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_937);
STATE_REG_938 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_938 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(938) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_938);
STATE_REG_939 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_939 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(939) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_939);
STATE_REG_940 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_940 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(940) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_940);
STATE_REG_941 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_941 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(941) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_941);
STATE_REG_942 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_942 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(942) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_942);
STATE_REG_943 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_943 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(943) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_943);
STATE_REG_944 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_944 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(944) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_944);
STATE_REG_945 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_945 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(945) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_945);
STATE_REG_946 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_946 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(946) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_946);
STATE_REG_947 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_947 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(947) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_947);
STATE_REG_948 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_948 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(948) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_948);
STATE_REG_949 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_949 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(949) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_949);
STATE_REG_950 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_950 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(950) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_950);
STATE_REG_951 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_951 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(951) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_951);
STATE_REG_952 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_952 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(952) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_952);
STATE_REG_953 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_953 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(953) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_953);
STATE_REG_954 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_954 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(954) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_954);
STATE_REG_955 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_955 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(955) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_955);
STATE_REG_956 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_956 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(956) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_956);
STATE_REG_957 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_957 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(957) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_957);
STATE_REG_958 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_958 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(958) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_958);
STATE_REG_959 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_959 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(959) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_959);
STATE_REG_960 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_960 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(960) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_960);
STATE_REG_961 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_961 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(961) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_961);
STATE_REG_962 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_962 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(962) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_962);
STATE_REG_963 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_963 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(963) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_963);
STATE_REG_964 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_964 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(964) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_964);
STATE_REG_965 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_965 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(965) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_965);
STATE_REG_966 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_966 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(966) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_966);
STATE_REG_967 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_967 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(967) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_967);
STATE_REG_968 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_968 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(968) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_968);
STATE_REG_969 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_969 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(969) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_969);
STATE_REG_970 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_970 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(970) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_970);
STATE_REG_971 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_971 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(971) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_971);
STATE_REG_972 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_972 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(972) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_972);
STATE_REG_973 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_973 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(973) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_973);
STATE_REG_974 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_974 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(974) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_974);
STATE_REG_975 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_975 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(975) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_975);
STATE_REG_976 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_976 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(976) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_976);
STATE_REG_977 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_977 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(977) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_977);
STATE_REG_978 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_978 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(978) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_978);
STATE_REG_979 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_979 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(979) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_979);
STATE_REG_980 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_980 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(980) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_980);
STATE_REG_981 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_981 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(981) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_981);
STATE_REG_982 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_982 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(982) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_982);
STATE_REG_983 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_983 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(983) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_983);
STATE_REG_984 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_984 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(984) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_984);
STATE_REG_985 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_985 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(985) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_985);
STATE_REG_986 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_986 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(986) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_986);
STATE_REG_987 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_987 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(987) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_987);
STATE_REG_988 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_988 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(988) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_988);
STATE_REG_989 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_989 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(989) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_989);
STATE_REG_990 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_990 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(990) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_990);
STATE_REG_991 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_991 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(991) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_991);
STATE_REG_992 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_992 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(992) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_992);
STATE_REG_993 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_993 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(993) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_993);
STATE_REG_994 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_994 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(994) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_994);
STATE_REG_995 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_995 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(995) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_995);
STATE_REG_996 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_996 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(996) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_996);
STATE_REG_997 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_997 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(997) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_997);
STATE_REG_998 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_998 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(998) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_998);
STATE_REG_999 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_999 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(999) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_999);
STATE_REG_1000 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1000 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1000) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1000);
STATE_REG_1001 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1001 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1001) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1001);
STATE_REG_1002 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1002 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1002) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1002);
STATE_REG_1003 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1003 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1003) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1003);
STATE_REG_1004 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1004 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1004) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1004);
STATE_REG_1005 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1005 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1005) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1005);
STATE_REG_1006 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1006 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1006) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1006);
STATE_REG_1007 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1007 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1007) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1007);
STATE_REG_1008 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1008 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1008) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1008);
STATE_REG_1009 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1009 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1009) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1009);
STATE_REG_1010 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1010 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1010) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1010);
STATE_REG_1011 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1011 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1011) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1011);
STATE_REG_1012 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1012 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1012) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1012);
STATE_REG_1013 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1013 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1013) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1013);
STATE_REG_1014 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1014 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1014) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1014);
STATE_REG_1015 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1015 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1015) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1015);
STATE_REG_1016 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1016 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1016) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1016);
STATE_REG_1017 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1017 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1017) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1017);
STATE_REG_1018 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1018 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1018) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1018);
STATE_REG_1019 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1019 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1019) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1019);
STATE_REG_1020 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1020 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1020) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1020);
STATE_REG_1021 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1021 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1021) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1021);
STATE_REG_1022 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1022 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1022) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1022);
STATE_REG_1023 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1023 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1023) ,
												REG_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1023);


MUX_SEL_UNIT_0 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_0 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_0 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_0
									);
MUX_SEL_UNIT_1 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_512 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1
									);
MUX_SEL_UNIT_2 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_2
									);
MUX_SEL_UNIT_3 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_513 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_3
									);
MUX_SEL_UNIT_4 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_2 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_2 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_4
									);
MUX_SEL_UNIT_5 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_514 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_5
									);
MUX_SEL_UNIT_6 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_3 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_3 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_6
									);
MUX_SEL_UNIT_7 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_515 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_7
									);
MUX_SEL_UNIT_8 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_4 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_4 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_8
									);
MUX_SEL_UNIT_9 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_516 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_9
									);
MUX_SEL_UNIT_10 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_5 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_5 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_10
									);
MUX_SEL_UNIT_11 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_517 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_11
									);
MUX_SEL_UNIT_12 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_6 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_6 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_12
									);
MUX_SEL_UNIT_13 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_518 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_13
									);
MUX_SEL_UNIT_14 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_7 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_7 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_14
									);
MUX_SEL_UNIT_15 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_519 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_15
									);
MUX_SEL_UNIT_16 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_8 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_8 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_16
									);
MUX_SEL_UNIT_17 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_520 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_17
									);
MUX_SEL_UNIT_18 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_9 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_9 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_18
									);
MUX_SEL_UNIT_19 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_521 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_19
									);
MUX_SEL_UNIT_20 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_10 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_10 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_20
									);
MUX_SEL_UNIT_21 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_522 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_21
									);
MUX_SEL_UNIT_22 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_11 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_11 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_22
									);
MUX_SEL_UNIT_23 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_523 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_23
									);
MUX_SEL_UNIT_24 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_12 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_12 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_24
									);
MUX_SEL_UNIT_25 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_524 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_25
									);
MUX_SEL_UNIT_26 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_13 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_13 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_26
									);
MUX_SEL_UNIT_27 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_525 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_27
									);
MUX_SEL_UNIT_28 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_14 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_14 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_28
									);
MUX_SEL_UNIT_29 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_526 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_29
									);
MUX_SEL_UNIT_30 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_15 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_15 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_30
									);
MUX_SEL_UNIT_31 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_527 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_31
									);
MUX_SEL_UNIT_32 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_16 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_16 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_32
									);
MUX_SEL_UNIT_33 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_528 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_33
									);
MUX_SEL_UNIT_34 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_17 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_17 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_34
									);
MUX_SEL_UNIT_35 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_529 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_35
									);
MUX_SEL_UNIT_36 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_18 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_18 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_36
									);
MUX_SEL_UNIT_37 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_530 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_37
									);
MUX_SEL_UNIT_38 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_19 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_19 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_38
									);
MUX_SEL_UNIT_39 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_531 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_39
									);
MUX_SEL_UNIT_40 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_20 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_20 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_40
									);
MUX_SEL_UNIT_41 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_532 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_41
									);
MUX_SEL_UNIT_42 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_21 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_21 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_42
									);
MUX_SEL_UNIT_43 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_533 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_43
									);
MUX_SEL_UNIT_44 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_22 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_22 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_44
									);
MUX_SEL_UNIT_45 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_534 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_45
									);
MUX_SEL_UNIT_46 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_23 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_23 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_46
									);
MUX_SEL_UNIT_47 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_535 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_47
									);
MUX_SEL_UNIT_48 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_24 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_24 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_48
									);
MUX_SEL_UNIT_49 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_536 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_49
									);
MUX_SEL_UNIT_50 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_25 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_25 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_50
									);
MUX_SEL_UNIT_51 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_537 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_51
									);
MUX_SEL_UNIT_52 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_26 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_26 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_52
									);
MUX_SEL_UNIT_53 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_538 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_53
									);
MUX_SEL_UNIT_54 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_27 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_27 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_54
									);
MUX_SEL_UNIT_55 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_539 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_55
									);
MUX_SEL_UNIT_56 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_28 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_28 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_56
									);
MUX_SEL_UNIT_57 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_540 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_57
									);
MUX_SEL_UNIT_58 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_29 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_29 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_58
									);
MUX_SEL_UNIT_59 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_541 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_59
									);
MUX_SEL_UNIT_60 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_30 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_30 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_60
									);
MUX_SEL_UNIT_61 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_542 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_61
									);
MUX_SEL_UNIT_62 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_31 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_31 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_62
									);
MUX_SEL_UNIT_63 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_543 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_63
									);
MUX_SEL_UNIT_64 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_32 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_32 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_64
									);
MUX_SEL_UNIT_65 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_544 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_65
									);
MUX_SEL_UNIT_66 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_33 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_33 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_66
									);
MUX_SEL_UNIT_67 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_545 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_67
									);
MUX_SEL_UNIT_68 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_34 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_34 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_68
									);
MUX_SEL_UNIT_69 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_546 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_69
									);
MUX_SEL_UNIT_70 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_35 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_35 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_70
									);
MUX_SEL_UNIT_71 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_547 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_71
									);
MUX_SEL_UNIT_72 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_36 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_36 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_72
									);
MUX_SEL_UNIT_73 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_548 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_73
									);
MUX_SEL_UNIT_74 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_37 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_37 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_74
									);
MUX_SEL_UNIT_75 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_549 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_75
									);
MUX_SEL_UNIT_76 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_38 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_38 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_76
									);
MUX_SEL_UNIT_77 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_550 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_77
									);
MUX_SEL_UNIT_78 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_39 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_39 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_78
									);
MUX_SEL_UNIT_79 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_551 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_79
									);
MUX_SEL_UNIT_80 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_40 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_40 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_80
									);
MUX_SEL_UNIT_81 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_552 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_81
									);
MUX_SEL_UNIT_82 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_41 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_41 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_82
									);
MUX_SEL_UNIT_83 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_553 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_83
									);
MUX_SEL_UNIT_84 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_42 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_42 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_84
									);
MUX_SEL_UNIT_85 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_554 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_85
									);
MUX_SEL_UNIT_86 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_43 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_43 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_86
									);
MUX_SEL_UNIT_87 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_555 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_87
									);
MUX_SEL_UNIT_88 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_44 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_44 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_88
									);
MUX_SEL_UNIT_89 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_556 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_89
									);
MUX_SEL_UNIT_90 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_45 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_45 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_90
									);
MUX_SEL_UNIT_91 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_557 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_91
									);
MUX_SEL_UNIT_92 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_46 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_46 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_92
									);
MUX_SEL_UNIT_93 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_558 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_93
									);
MUX_SEL_UNIT_94 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_47 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_47 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_94
									);
MUX_SEL_UNIT_95 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_559 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_95
									);
MUX_SEL_UNIT_96 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_48 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_48 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_96
									);
MUX_SEL_UNIT_97 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_560 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_97
									);
MUX_SEL_UNIT_98 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_49 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_49 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_98
									);
MUX_SEL_UNIT_99 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_561 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_99
									);
MUX_SEL_UNIT_100 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_50 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_50 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_100
									);
MUX_SEL_UNIT_101 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_562 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_101
									);
MUX_SEL_UNIT_102 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_51 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_51 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_102
									);
MUX_SEL_UNIT_103 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_563 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_103
									);
MUX_SEL_UNIT_104 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_52 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_52 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_104
									);
MUX_SEL_UNIT_105 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_564 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_105
									);
MUX_SEL_UNIT_106 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_53 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_53 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_106
									);
MUX_SEL_UNIT_107 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_565 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_107
									);
MUX_SEL_UNIT_108 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_54 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_54 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_108
									);
MUX_SEL_UNIT_109 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_566 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_109
									);
MUX_SEL_UNIT_110 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_55 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_55 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_110
									);
MUX_SEL_UNIT_111 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_567 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_111
									);
MUX_SEL_UNIT_112 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_56 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_56 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_112
									);
MUX_SEL_UNIT_113 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_568 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_113
									);
MUX_SEL_UNIT_114 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_57 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_57 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_114
									);
MUX_SEL_UNIT_115 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_569 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_115
									);
MUX_SEL_UNIT_116 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_58 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_58 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_116
									);
MUX_SEL_UNIT_117 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_570 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_117
									);
MUX_SEL_UNIT_118 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_59 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_59 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_118
									);
MUX_SEL_UNIT_119 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_571 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_119
									);
MUX_SEL_UNIT_120 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_60 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_60 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_120
									);
MUX_SEL_UNIT_121 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_572 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_121
									);
MUX_SEL_UNIT_122 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_61 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_61 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_122
									);
MUX_SEL_UNIT_123 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_573 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_123
									);
MUX_SEL_UNIT_124 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_62 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_62 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_124
									);
MUX_SEL_UNIT_125 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_574 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_125
									);
MUX_SEL_UNIT_126 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_63 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_63 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_126
									);
MUX_SEL_UNIT_127 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_575 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_127
									);
MUX_SEL_UNIT_128 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_64 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_64 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_128
									);
MUX_SEL_UNIT_129 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_576 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_129
									);
MUX_SEL_UNIT_130 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_65 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_65 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_130
									);
MUX_SEL_UNIT_131 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_577 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_131
									);
MUX_SEL_UNIT_132 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_66 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_66 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_132
									);
MUX_SEL_UNIT_133 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_578 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_133
									);
MUX_SEL_UNIT_134 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_67 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_67 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_134
									);
MUX_SEL_UNIT_135 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_579 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_135
									);
MUX_SEL_UNIT_136 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_68 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_68 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_136
									);
MUX_SEL_UNIT_137 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_580 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_137
									);
MUX_SEL_UNIT_138 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_69 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_69 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_138
									);
MUX_SEL_UNIT_139 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_581 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_139
									);
MUX_SEL_UNIT_140 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_70 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_70 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_140
									);
MUX_SEL_UNIT_141 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_582 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_141
									);
MUX_SEL_UNIT_142 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_71 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_71 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_142
									);
MUX_SEL_UNIT_143 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_583 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_143
									);
MUX_SEL_UNIT_144 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_72 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_72 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_144
									);
MUX_SEL_UNIT_145 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_584 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_145
									);
MUX_SEL_UNIT_146 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_73 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_73 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_146
									);
MUX_SEL_UNIT_147 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_585 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_147
									);
MUX_SEL_UNIT_148 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_74 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_74 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_148
									);
MUX_SEL_UNIT_149 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_586 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_149
									);
MUX_SEL_UNIT_150 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_75 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_75 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_150
									);
MUX_SEL_UNIT_151 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_587 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_151
									);
MUX_SEL_UNIT_152 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_76 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_76 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_152
									);
MUX_SEL_UNIT_153 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_588 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_153
									);
MUX_SEL_UNIT_154 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_77 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_77 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_154
									);
MUX_SEL_UNIT_155 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_589 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_155
									);
MUX_SEL_UNIT_156 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_78 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_78 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_156
									);
MUX_SEL_UNIT_157 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_590 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_157
									);
MUX_SEL_UNIT_158 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_79 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_79 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_158
									);
MUX_SEL_UNIT_159 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_591 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_159
									);
MUX_SEL_UNIT_160 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_80 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_80 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_160
									);
MUX_SEL_UNIT_161 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_592 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_161
									);
MUX_SEL_UNIT_162 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_81 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_81 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_162
									);
MUX_SEL_UNIT_163 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_593 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_163
									);
MUX_SEL_UNIT_164 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_82 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_82 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_164
									);
MUX_SEL_UNIT_165 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_594 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_165
									);
MUX_SEL_UNIT_166 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_83 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_83 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_166
									);
MUX_SEL_UNIT_167 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_595 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_167
									);
MUX_SEL_UNIT_168 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_84 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_84 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_168
									);
MUX_SEL_UNIT_169 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_596 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_169
									);
MUX_SEL_UNIT_170 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_85 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_85 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_170
									);
MUX_SEL_UNIT_171 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_597 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_171
									);
MUX_SEL_UNIT_172 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_86 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_86 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_172
									);
MUX_SEL_UNIT_173 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_598 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_173
									);
MUX_SEL_UNIT_174 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_87 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_87 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_174
									);
MUX_SEL_UNIT_175 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_599 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_175
									);
MUX_SEL_UNIT_176 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_88 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_88 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_176
									);
MUX_SEL_UNIT_177 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_600 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_177
									);
MUX_SEL_UNIT_178 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_89 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_89 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_178
									);
MUX_SEL_UNIT_179 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_601 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_179
									);
MUX_SEL_UNIT_180 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_90 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_90 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_180
									);
MUX_SEL_UNIT_181 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_602 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_181
									);
MUX_SEL_UNIT_182 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_91 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_91 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_182
									);
MUX_SEL_UNIT_183 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_603 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_183
									);
MUX_SEL_UNIT_184 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_92 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_92 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_184
									);
MUX_SEL_UNIT_185 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_604 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_185
									);
MUX_SEL_UNIT_186 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_93 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_93 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_186
									);
MUX_SEL_UNIT_187 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_605 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_187
									);
MUX_SEL_UNIT_188 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_94 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_94 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_188
									);
MUX_SEL_UNIT_189 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_606 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_189
									);
MUX_SEL_UNIT_190 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_95 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_95 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_190
									);
MUX_SEL_UNIT_191 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_607 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_191
									);
MUX_SEL_UNIT_192 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_96 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_96 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_192
									);
MUX_SEL_UNIT_193 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_608 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_193
									);
MUX_SEL_UNIT_194 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_97 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_97 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_194
									);
MUX_SEL_UNIT_195 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_609 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_195
									);
MUX_SEL_UNIT_196 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_98 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_98 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_196
									);
MUX_SEL_UNIT_197 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_610 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_197
									);
MUX_SEL_UNIT_198 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_99 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_99 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_198
									);
MUX_SEL_UNIT_199 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_611 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_199
									);
MUX_SEL_UNIT_200 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_100 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_100 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_200
									);
MUX_SEL_UNIT_201 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_612 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_201
									);
MUX_SEL_UNIT_202 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_101 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_101 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_202
									);
MUX_SEL_UNIT_203 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_613 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_203
									);
MUX_SEL_UNIT_204 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_102 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_102 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_204
									);
MUX_SEL_UNIT_205 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_614 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_205
									);
MUX_SEL_UNIT_206 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_103 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_103 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_206
									);
MUX_SEL_UNIT_207 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_615 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_207
									);
MUX_SEL_UNIT_208 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_104 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_104 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_208
									);
MUX_SEL_UNIT_209 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_616 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_209
									);
MUX_SEL_UNIT_210 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_105 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_105 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_210
									);
MUX_SEL_UNIT_211 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_617 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_211
									);
MUX_SEL_UNIT_212 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_106 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_106 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_212
									);
MUX_SEL_UNIT_213 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_618 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_213
									);
MUX_SEL_UNIT_214 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_107 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_107 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_214
									);
MUX_SEL_UNIT_215 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_619 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_215
									);
MUX_SEL_UNIT_216 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_108 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_108 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_216
									);
MUX_SEL_UNIT_217 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_620 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_217
									);
MUX_SEL_UNIT_218 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_109 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_109 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_218
									);
MUX_SEL_UNIT_219 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_621 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_219
									);
MUX_SEL_UNIT_220 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_110 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_110 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_220
									);
MUX_SEL_UNIT_221 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_622 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_221
									);
MUX_SEL_UNIT_222 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_111 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_111 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_222
									);
MUX_SEL_UNIT_223 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_623 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_223
									);
MUX_SEL_UNIT_224 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_112 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_112 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_224
									);
MUX_SEL_UNIT_225 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_624 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_225
									);
MUX_SEL_UNIT_226 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_113 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_113 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_226
									);
MUX_SEL_UNIT_227 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_625 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_227
									);
MUX_SEL_UNIT_228 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_114 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_114 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_228
									);
MUX_SEL_UNIT_229 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_626 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_229
									);
MUX_SEL_UNIT_230 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_115 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_115 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_230
									);
MUX_SEL_UNIT_231 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_627 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_231
									);
MUX_SEL_UNIT_232 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_116 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_116 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_232
									);
MUX_SEL_UNIT_233 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_628 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_233
									);
MUX_SEL_UNIT_234 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_117 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_117 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_234
									);
MUX_SEL_UNIT_235 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_629 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_235
									);
MUX_SEL_UNIT_236 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_118 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_118 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_236
									);
MUX_SEL_UNIT_237 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_630 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_237
									);
MUX_SEL_UNIT_238 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_119 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_119 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_238
									);
MUX_SEL_UNIT_239 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_631 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_239
									);
MUX_SEL_UNIT_240 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_120 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_120 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_240
									);
MUX_SEL_UNIT_241 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_632 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_241
									);
MUX_SEL_UNIT_242 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_121 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_121 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_242
									);
MUX_SEL_UNIT_243 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_633 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_243
									);
MUX_SEL_UNIT_244 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_122 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_122 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_244
									);
MUX_SEL_UNIT_245 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_634 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_245
									);
MUX_SEL_UNIT_246 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_123 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_123 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_246
									);
MUX_SEL_UNIT_247 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_635 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_247
									);
MUX_SEL_UNIT_248 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_124 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_124 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_248
									);
MUX_SEL_UNIT_249 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_636 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_249
									);
MUX_SEL_UNIT_250 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_125 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_125 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_250
									);
MUX_SEL_UNIT_251 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_637 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_251
									);
MUX_SEL_UNIT_252 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_126 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_126 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_252
									);
MUX_SEL_UNIT_253 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_638 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_253
									);
MUX_SEL_UNIT_254 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_127 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_127 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_254
									);
MUX_SEL_UNIT_255 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_639 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_255
									);
MUX_SEL_UNIT_256 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_256 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_128 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_128 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_256
									);
MUX_SEL_UNIT_257 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_640 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_257
									);
MUX_SEL_UNIT_258 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_257 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_129 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_129 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_258
									);
MUX_SEL_UNIT_259 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_641 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_259
									);
MUX_SEL_UNIT_260 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_258 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_130 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_130 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_260
									);
MUX_SEL_UNIT_261 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_642 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_261
									);
MUX_SEL_UNIT_262 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_259 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_131 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_131 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_262
									);
MUX_SEL_UNIT_263 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_643 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_263
									);
MUX_SEL_UNIT_264 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_260 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_132 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_132 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_264
									);
MUX_SEL_UNIT_265 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_644 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_265
									);
MUX_SEL_UNIT_266 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_261 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_133 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_133 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_266
									);
MUX_SEL_UNIT_267 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_645 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_267
									);
MUX_SEL_UNIT_268 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_262 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_134 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_134 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_268
									);
MUX_SEL_UNIT_269 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_646 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_269
									);
MUX_SEL_UNIT_270 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_263 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_135 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_135 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_270
									);
MUX_SEL_UNIT_271 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_647 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_271
									);
MUX_SEL_UNIT_272 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_264 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_136 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_136 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_272
									);
MUX_SEL_UNIT_273 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_648 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_273
									);
MUX_SEL_UNIT_274 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_265 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_137 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_137 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_274
									);
MUX_SEL_UNIT_275 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_649 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_275
									);
MUX_SEL_UNIT_276 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_266 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_138 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_138 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_276
									);
MUX_SEL_UNIT_277 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_650 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_277
									);
MUX_SEL_UNIT_278 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_267 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_139 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_139 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_278
									);
MUX_SEL_UNIT_279 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_651 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_279
									);
MUX_SEL_UNIT_280 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_268 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_140 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_140 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_280
									);
MUX_SEL_UNIT_281 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_652 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_281
									);
MUX_SEL_UNIT_282 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_269 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_141 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_141 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_282
									);
MUX_SEL_UNIT_283 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_653 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_283
									);
MUX_SEL_UNIT_284 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_270 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_142 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_142 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_284
									);
MUX_SEL_UNIT_285 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_654 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_285
									);
MUX_SEL_UNIT_286 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_271 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_143 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_143 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_286
									);
MUX_SEL_UNIT_287 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_655 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_287
									);
MUX_SEL_UNIT_288 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_272 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_144 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_144 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_288
									);
MUX_SEL_UNIT_289 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_656 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_289
									);
MUX_SEL_UNIT_290 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_273 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_145 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_145 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_290
									);
MUX_SEL_UNIT_291 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_657 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_291
									);
MUX_SEL_UNIT_292 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_274 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_146 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_146 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_292
									);
MUX_SEL_UNIT_293 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_658 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_293
									);
MUX_SEL_UNIT_294 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_275 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_147 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_147 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_294
									);
MUX_SEL_UNIT_295 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_659 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_295
									);
MUX_SEL_UNIT_296 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_276 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_148 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_148 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_296
									);
MUX_SEL_UNIT_297 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_660 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_297
									);
MUX_SEL_UNIT_298 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_277 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_149 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_149 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_298
									);
MUX_SEL_UNIT_299 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_661 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_299
									);
MUX_SEL_UNIT_300 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_278 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_150 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_150 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_300
									);
MUX_SEL_UNIT_301 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_662 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_301
									);
MUX_SEL_UNIT_302 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_279 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_151 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_151 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_302
									);
MUX_SEL_UNIT_303 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_663 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_303
									);
MUX_SEL_UNIT_304 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_280 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_152 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_152 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_304
									);
MUX_SEL_UNIT_305 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_664 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_305
									);
MUX_SEL_UNIT_306 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_281 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_153 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_153 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_306
									);
MUX_SEL_UNIT_307 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_665 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_307
									);
MUX_SEL_UNIT_308 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_282 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_154 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_154 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_308
									);
MUX_SEL_UNIT_309 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_666 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_309
									);
MUX_SEL_UNIT_310 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_283 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_155 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_155 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_310
									);
MUX_SEL_UNIT_311 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_667 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_311
									);
MUX_SEL_UNIT_312 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_284 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_156 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_156 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_312
									);
MUX_SEL_UNIT_313 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_668 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_313
									);
MUX_SEL_UNIT_314 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_285 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_157 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_157 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_314
									);
MUX_SEL_UNIT_315 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_669 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_315
									);
MUX_SEL_UNIT_316 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_286 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_158 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_158 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_316
									);
MUX_SEL_UNIT_317 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_670 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_317
									);
MUX_SEL_UNIT_318 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_287 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_159 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_159 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_318
									);
MUX_SEL_UNIT_319 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_671 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_319
									);
MUX_SEL_UNIT_320 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_288 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_160 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_160 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_320
									);
MUX_SEL_UNIT_321 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_672 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_321
									);
MUX_SEL_UNIT_322 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_289 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_161 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_161 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_322
									);
MUX_SEL_UNIT_323 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_673 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_323
									);
MUX_SEL_UNIT_324 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_290 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_162 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_162 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_324
									);
MUX_SEL_UNIT_325 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_674 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_325
									);
MUX_SEL_UNIT_326 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_291 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_163 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_163 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_326
									);
MUX_SEL_UNIT_327 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_675 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_327
									);
MUX_SEL_UNIT_328 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_292 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_164 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_164 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_328
									);
MUX_SEL_UNIT_329 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_676 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_329
									);
MUX_SEL_UNIT_330 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_293 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_165 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_165 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_330
									);
MUX_SEL_UNIT_331 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_677 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_331
									);
MUX_SEL_UNIT_332 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_294 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_166 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_166 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_332
									);
MUX_SEL_UNIT_333 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_678 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_333
									);
MUX_SEL_UNIT_334 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_295 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_167 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_167 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_334
									);
MUX_SEL_UNIT_335 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_679 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_335
									);
MUX_SEL_UNIT_336 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_296 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_168 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_168 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_336
									);
MUX_SEL_UNIT_337 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_680 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_337
									);
MUX_SEL_UNIT_338 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_297 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_169 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_169 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_338
									);
MUX_SEL_UNIT_339 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_681 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_339
									);
MUX_SEL_UNIT_340 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_298 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_170 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_170 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_340
									);
MUX_SEL_UNIT_341 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_682 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_341
									);
MUX_SEL_UNIT_342 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_299 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_171 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_171 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_342
									);
MUX_SEL_UNIT_343 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_683 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_343
									);
MUX_SEL_UNIT_344 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_300 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_172 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_172 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_344
									);
MUX_SEL_UNIT_345 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_684 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_345
									);
MUX_SEL_UNIT_346 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_301 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_173 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_173 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_346
									);
MUX_SEL_UNIT_347 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_685 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_347
									);
MUX_SEL_UNIT_348 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_302 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_174 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_174 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_348
									);
MUX_SEL_UNIT_349 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_686 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_349
									);
MUX_SEL_UNIT_350 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_303 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_175 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_175 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_350
									);
MUX_SEL_UNIT_351 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_687 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_351
									);
MUX_SEL_UNIT_352 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_304 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_176 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_176 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_352
									);
MUX_SEL_UNIT_353 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_688 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_353
									);
MUX_SEL_UNIT_354 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_305 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_177 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_177 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_354
									);
MUX_SEL_UNIT_355 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_689 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_355
									);
MUX_SEL_UNIT_356 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_306 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_178 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_178 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_356
									);
MUX_SEL_UNIT_357 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_690 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_357
									);
MUX_SEL_UNIT_358 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_307 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_179 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_179 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_358
									);
MUX_SEL_UNIT_359 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_691 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_359
									);
MUX_SEL_UNIT_360 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_308 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_180 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_180 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_360
									);
MUX_SEL_UNIT_361 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_692 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_361
									);
MUX_SEL_UNIT_362 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_309 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_181 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_181 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_362
									);
MUX_SEL_UNIT_363 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_693 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_363
									);
MUX_SEL_UNIT_364 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_310 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_182 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_182 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_364
									);
MUX_SEL_UNIT_365 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_694 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_365
									);
MUX_SEL_UNIT_366 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_311 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_183 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_183 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_366
									);
MUX_SEL_UNIT_367 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_695 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_367
									);
MUX_SEL_UNIT_368 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_312 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_184 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_184 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_368
									);
MUX_SEL_UNIT_369 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_696 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_369
									);
MUX_SEL_UNIT_370 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_313 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_185 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_185 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_370
									);
MUX_SEL_UNIT_371 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_697 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_371
									);
MUX_SEL_UNIT_372 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_314 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_186 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_186 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_372
									);
MUX_SEL_UNIT_373 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_698 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_373
									);
MUX_SEL_UNIT_374 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_315 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_187 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_187 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_374
									);
MUX_SEL_UNIT_375 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_699 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_375
									);
MUX_SEL_UNIT_376 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_316 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_188 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_188 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_376
									);
MUX_SEL_UNIT_377 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_700 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_377
									);
MUX_SEL_UNIT_378 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_317 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_189 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_189 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_378
									);
MUX_SEL_UNIT_379 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_701 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_379
									);
MUX_SEL_UNIT_380 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_318 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_190 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_190 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_380
									);
MUX_SEL_UNIT_381 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_702 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_381
									);
MUX_SEL_UNIT_382 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_319 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_191 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_191 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_382
									);
MUX_SEL_UNIT_383 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_703 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_383
									);
MUX_SEL_UNIT_384 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_384 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_320 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_192 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_192 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_384
									);
MUX_SEL_UNIT_385 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_704 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_385
									);
MUX_SEL_UNIT_386 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_385 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_321 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_193 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_193 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_386
									);
MUX_SEL_UNIT_387 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_705 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_387
									);
MUX_SEL_UNIT_388 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_386 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_322 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_194 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_194 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_388
									);
MUX_SEL_UNIT_389 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_706 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_389
									);
MUX_SEL_UNIT_390 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_387 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_323 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_195 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_195 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_390
									);
MUX_SEL_UNIT_391 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_707 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_391
									);
MUX_SEL_UNIT_392 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_388 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_324 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_196 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_196 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_392
									);
MUX_SEL_UNIT_393 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_708 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_393
									);
MUX_SEL_UNIT_394 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_389 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_325 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_197 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_197 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_394
									);
MUX_SEL_UNIT_395 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_709 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_395
									);
MUX_SEL_UNIT_396 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_390 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_326 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_198 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_198 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_396
									);
MUX_SEL_UNIT_397 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_710 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_397
									);
MUX_SEL_UNIT_398 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_391 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_327 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_199 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_199 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_398
									);
MUX_SEL_UNIT_399 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_711 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_399
									);
MUX_SEL_UNIT_400 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_392 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_328 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_200 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_200 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_400
									);
MUX_SEL_UNIT_401 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_712 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_401
									);
MUX_SEL_UNIT_402 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_393 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_329 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_201 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_201 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_402
									);
MUX_SEL_UNIT_403 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_713 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_403
									);
MUX_SEL_UNIT_404 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_394 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_330 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_202 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_202 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_404
									);
MUX_SEL_UNIT_405 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_714 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_405
									);
MUX_SEL_UNIT_406 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_395 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_331 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_203 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_203 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_406
									);
MUX_SEL_UNIT_407 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_715 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_407
									);
MUX_SEL_UNIT_408 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_396 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_332 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_204 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_204 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_408
									);
MUX_SEL_UNIT_409 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_716 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_409
									);
MUX_SEL_UNIT_410 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_397 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_333 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_205 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_205 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_410
									);
MUX_SEL_UNIT_411 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_717 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_411
									);
MUX_SEL_UNIT_412 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_398 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_334 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_206 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_206 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_412
									);
MUX_SEL_UNIT_413 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_718 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_413
									);
MUX_SEL_UNIT_414 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_399 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_335 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_207 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_207 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_414
									);
MUX_SEL_UNIT_415 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_719 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_415
									);
MUX_SEL_UNIT_416 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_400 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_336 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_208 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_208 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_416
									);
MUX_SEL_UNIT_417 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_720 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_417
									);
MUX_SEL_UNIT_418 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_401 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_337 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_209 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_209 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_418
									);
MUX_SEL_UNIT_419 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_721 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_419
									);
MUX_SEL_UNIT_420 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_402 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_338 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_210 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_210 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_420
									);
MUX_SEL_UNIT_421 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_722 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_421
									);
MUX_SEL_UNIT_422 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_403 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_339 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_211 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_211 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_422
									);
MUX_SEL_UNIT_423 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_723 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_423
									);
MUX_SEL_UNIT_424 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_404 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_340 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_212 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_212 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_424
									);
MUX_SEL_UNIT_425 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_724 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_425
									);
MUX_SEL_UNIT_426 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_405 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_341 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_213 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_213 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_426
									);
MUX_SEL_UNIT_427 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_725 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_427
									);
MUX_SEL_UNIT_428 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_406 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_342 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_214 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_214 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_428
									);
MUX_SEL_UNIT_429 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_726 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_429
									);
MUX_SEL_UNIT_430 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_407 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_343 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_215 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_215 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_430
									);
MUX_SEL_UNIT_431 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_727 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_431
									);
MUX_SEL_UNIT_432 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_408 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_344 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_216 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_216 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_432
									);
MUX_SEL_UNIT_433 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_728 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_433
									);
MUX_SEL_UNIT_434 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_409 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_345 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_217 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_217 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_434
									);
MUX_SEL_UNIT_435 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_729 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_435
									);
MUX_SEL_UNIT_436 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_410 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_346 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_218 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_218 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_436
									);
MUX_SEL_UNIT_437 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_730 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_437
									);
MUX_SEL_UNIT_438 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_411 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_347 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_219 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_219 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_438
									);
MUX_SEL_UNIT_439 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_731 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_439
									);
MUX_SEL_UNIT_440 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_412 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_348 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_220 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_220 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_440
									);
MUX_SEL_UNIT_441 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_732 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_441
									);
MUX_SEL_UNIT_442 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_413 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_349 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_221 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_221 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_442
									);
MUX_SEL_UNIT_443 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_733 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_443
									);
MUX_SEL_UNIT_444 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_414 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_350 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_222 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_222 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_444
									);
MUX_SEL_UNIT_445 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_734 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_445
									);
MUX_SEL_UNIT_446 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_415 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_351 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_223 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_223 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_446
									);
MUX_SEL_UNIT_447 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_735 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_447
									);
MUX_SEL_UNIT_448 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_448 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_416 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_352 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_224 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_224 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_448
									);
MUX_SEL_UNIT_449 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_736 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_449
									);
MUX_SEL_UNIT_450 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_449 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_417 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_353 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_225 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_225 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_450
									);
MUX_SEL_UNIT_451 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_737 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_451
									);
MUX_SEL_UNIT_452 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_450 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_418 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_354 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_226 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_226 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_452
									);
MUX_SEL_UNIT_453 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_738 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_453
									);
MUX_SEL_UNIT_454 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_451 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_419 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_355 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_227 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_227 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_454
									);
MUX_SEL_UNIT_455 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_739 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_455
									);
MUX_SEL_UNIT_456 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_452 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_420 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_356 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_228 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_228 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_456
									);
MUX_SEL_UNIT_457 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_740 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_457
									);
MUX_SEL_UNIT_458 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_453 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_421 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_357 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_229 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_229 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_458
									);
MUX_SEL_UNIT_459 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_741 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_459
									);
MUX_SEL_UNIT_460 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_454 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_422 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_358 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_230 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_230 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_460
									);
MUX_SEL_UNIT_461 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_742 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_461
									);
MUX_SEL_UNIT_462 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_455 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_423 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_359 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_231 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_231 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_462
									);
MUX_SEL_UNIT_463 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_743 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_463
									);
MUX_SEL_UNIT_464 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_456 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_424 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_360 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_232 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_232 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_464
									);
MUX_SEL_UNIT_465 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_744 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_465
									);
MUX_SEL_UNIT_466 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_457 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_425 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_361 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_233 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_233 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_466
									);
MUX_SEL_UNIT_467 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_745 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_467
									);
MUX_SEL_UNIT_468 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_458 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_426 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_362 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_234 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_234 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_468
									);
MUX_SEL_UNIT_469 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_746 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_469
									);
MUX_SEL_UNIT_470 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_459 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_427 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_363 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_235 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_235 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_470
									);
MUX_SEL_UNIT_471 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_747 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_471
									);
MUX_SEL_UNIT_472 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_460 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_428 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_364 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_236 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_236 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_472
									);
MUX_SEL_UNIT_473 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_748 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_473
									);
MUX_SEL_UNIT_474 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_461 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_429 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_365 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_237 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_237 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_474
									);
MUX_SEL_UNIT_475 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_749 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_475
									);
MUX_SEL_UNIT_476 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_462 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_430 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_366 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_238 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_238 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_476
									);
MUX_SEL_UNIT_477 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_750 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_477
									);
MUX_SEL_UNIT_478 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_463 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_431 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_367 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_239 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_239 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_478
									);
MUX_SEL_UNIT_479 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_751 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_479
									);
MUX_SEL_UNIT_480 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_480 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_464 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_432 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_368 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_240 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_240 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_480
									);
MUX_SEL_UNIT_481 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_752 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_481
									);
MUX_SEL_UNIT_482 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_481 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_465 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_433 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_369 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_241 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_241 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_482
									);
MUX_SEL_UNIT_483 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_753 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_483
									);
MUX_SEL_UNIT_484 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_482 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_466 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_434 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_370 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_242 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_242 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_484
									);
MUX_SEL_UNIT_485 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_754 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_485
									);
MUX_SEL_UNIT_486 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_483 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_467 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_435 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_371 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_243 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_243 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_486
									);
MUX_SEL_UNIT_487 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_755 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_487
									);
MUX_SEL_UNIT_488 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_484 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_468 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_436 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_372 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_244 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_244 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_488
									);
MUX_SEL_UNIT_489 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_756 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_489
									);
MUX_SEL_UNIT_490 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_485 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_469 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_437 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_373 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_245 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_245 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_490
									);
MUX_SEL_UNIT_491 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_757 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_491
									);
MUX_SEL_UNIT_492 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_486 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_470 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_438 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_374 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_246 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_246 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_492
									);
MUX_SEL_UNIT_493 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_758 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_493
									);
MUX_SEL_UNIT_494 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_487 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_471 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_439 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_375 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_247 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_247 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_494
									);
MUX_SEL_UNIT_495 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_759 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_495
									);
MUX_SEL_UNIT_496 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_496 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_488 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_472 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_440 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_376 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_248 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_248 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_496
									);
MUX_SEL_UNIT_497 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_760 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_497
									);
MUX_SEL_UNIT_498 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_497 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_489 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_473 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_441 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_377 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_249 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_249 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_498
									);
MUX_SEL_UNIT_499 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_761 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_499
									);
MUX_SEL_UNIT_500 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_498 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_490 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_474 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_442 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_378 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_250 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_250 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_500
									);
MUX_SEL_UNIT_501 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_762 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_501
									);
MUX_SEL_UNIT_502 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_499 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_491 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_475 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_443 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_379 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_251 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_251 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_502
									);
MUX_SEL_UNIT_503 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_763 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_503
									);
MUX_SEL_UNIT_504 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_504 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_500 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_492 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_476 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_444 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_380 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_252 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_252 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_504
									);
MUX_SEL_UNIT_505 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_764 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_505
									);
MUX_SEL_UNIT_506 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_505 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_501 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_493 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_477 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_445 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_381 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_253 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_253 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_506
									);
MUX_SEL_UNIT_507 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_765 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_507
									);
MUX_SEL_UNIT_508 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_508 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_506 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_502 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_494 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_478 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_446 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_382 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_254 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_254 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_508
									);
MUX_SEL_UNIT_509 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_766 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_509
									);
MUX_SEL_UNIT_510 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_510 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_509 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_507 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_503 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_495 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_479 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_447 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_383 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_255 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_255 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_510
									);
MUX_SEL_UNIT_511 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_511 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_767 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_511
									);
MUX_SEL_UNIT_512 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_512 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_256 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_512
									);
MUX_SEL_UNIT_513 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_768 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_513
									);
MUX_SEL_UNIT_514 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_513 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_257 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_514
									);
MUX_SEL_UNIT_515 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_769 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_515
									);
MUX_SEL_UNIT_516 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_514 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_258 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_516
									);
MUX_SEL_UNIT_517 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_770 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_517
									);
MUX_SEL_UNIT_518 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_515 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_259 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_518
									);
MUX_SEL_UNIT_519 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_771 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_519
									);
MUX_SEL_UNIT_520 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_516 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_260 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_520
									);
MUX_SEL_UNIT_521 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_772 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_521
									);
MUX_SEL_UNIT_522 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_517 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_261 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_522
									);
MUX_SEL_UNIT_523 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_773 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_523
									);
MUX_SEL_UNIT_524 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_518 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_262 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_524
									);
MUX_SEL_UNIT_525 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_774 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_525
									);
MUX_SEL_UNIT_526 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_519 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_263 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_526
									);
MUX_SEL_UNIT_527 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_775 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_527
									);
MUX_SEL_UNIT_528 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_520 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_264 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_528
									);
MUX_SEL_UNIT_529 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_776 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_529
									);
MUX_SEL_UNIT_530 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_521 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_265 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_530
									);
MUX_SEL_UNIT_531 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_777 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_531
									);
MUX_SEL_UNIT_532 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_522 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_266 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_532
									);
MUX_SEL_UNIT_533 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_778 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_533
									);
MUX_SEL_UNIT_534 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_523 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_267 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_534
									);
MUX_SEL_UNIT_535 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_779 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_535
									);
MUX_SEL_UNIT_536 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_524 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_268 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_536
									);
MUX_SEL_UNIT_537 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_780 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_537
									);
MUX_SEL_UNIT_538 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_525 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_269 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_538
									);
MUX_SEL_UNIT_539 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_781 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_539
									);
MUX_SEL_UNIT_540 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_526 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_270 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_540
									);
MUX_SEL_UNIT_541 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_782 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_541
									);
MUX_SEL_UNIT_542 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_527 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_271 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_542
									);
MUX_SEL_UNIT_543 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_783 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_543
									);
MUX_SEL_UNIT_544 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_528 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_272 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_544
									);
MUX_SEL_UNIT_545 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_784 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_545
									);
MUX_SEL_UNIT_546 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_529 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_273 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_546
									);
MUX_SEL_UNIT_547 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_785 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_547
									);
MUX_SEL_UNIT_548 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_530 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_274 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_548
									);
MUX_SEL_UNIT_549 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_786 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_549
									);
MUX_SEL_UNIT_550 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_531 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_275 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_550
									);
MUX_SEL_UNIT_551 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_787 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_551
									);
MUX_SEL_UNIT_552 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_532 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_276 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_552
									);
MUX_SEL_UNIT_553 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_788 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_553
									);
MUX_SEL_UNIT_554 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_533 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_277 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_554
									);
MUX_SEL_UNIT_555 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_789 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_555
									);
MUX_SEL_UNIT_556 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_534 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_278 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_556
									);
MUX_SEL_UNIT_557 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_790 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_557
									);
MUX_SEL_UNIT_558 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_535 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_279 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_558
									);
MUX_SEL_UNIT_559 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_791 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_559
									);
MUX_SEL_UNIT_560 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_536 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_280 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_560
									);
MUX_SEL_UNIT_561 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_792 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_561
									);
MUX_SEL_UNIT_562 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_537 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_281 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_562
									);
MUX_SEL_UNIT_563 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_793 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_563
									);
MUX_SEL_UNIT_564 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_538 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_282 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_564
									);
MUX_SEL_UNIT_565 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_794 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_565
									);
MUX_SEL_UNIT_566 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_539 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_283 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_566
									);
MUX_SEL_UNIT_567 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_795 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_567
									);
MUX_SEL_UNIT_568 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_540 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_284 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_568
									);
MUX_SEL_UNIT_569 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_796 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_569
									);
MUX_SEL_UNIT_570 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_541 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_285 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_570
									);
MUX_SEL_UNIT_571 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_797 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_571
									);
MUX_SEL_UNIT_572 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_542 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_286 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_572
									);
MUX_SEL_UNIT_573 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_798 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_573
									);
MUX_SEL_UNIT_574 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_543 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_287 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_574
									);
MUX_SEL_UNIT_575 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_799 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_575
									);
MUX_SEL_UNIT_576 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_544 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_288 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_576
									);
MUX_SEL_UNIT_577 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_800 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_577
									);
MUX_SEL_UNIT_578 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_545 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_289 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_578
									);
MUX_SEL_UNIT_579 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_801 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_579
									);
MUX_SEL_UNIT_580 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_546 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_290 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_580
									);
MUX_SEL_UNIT_581 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_802 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_581
									);
MUX_SEL_UNIT_582 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_547 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_291 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_582
									);
MUX_SEL_UNIT_583 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_803 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_583
									);
MUX_SEL_UNIT_584 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_548 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_292 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_584
									);
MUX_SEL_UNIT_585 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_804 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_585
									);
MUX_SEL_UNIT_586 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_549 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_293 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_586
									);
MUX_SEL_UNIT_587 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_805 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_587
									);
MUX_SEL_UNIT_588 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_550 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_294 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_588
									);
MUX_SEL_UNIT_589 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_806 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_589
									);
MUX_SEL_UNIT_590 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_551 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_295 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_590
									);
MUX_SEL_UNIT_591 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_807 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_591
									);
MUX_SEL_UNIT_592 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_552 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_296 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_592
									);
MUX_SEL_UNIT_593 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_808 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_593
									);
MUX_SEL_UNIT_594 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_553 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_297 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_594
									);
MUX_SEL_UNIT_595 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_809 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_595
									);
MUX_SEL_UNIT_596 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_554 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_298 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_596
									);
MUX_SEL_UNIT_597 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_810 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_597
									);
MUX_SEL_UNIT_598 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_555 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_299 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_598
									);
MUX_SEL_UNIT_599 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_811 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_599
									);
MUX_SEL_UNIT_600 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_556 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_300 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_600
									);
MUX_SEL_UNIT_601 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_812 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_601
									);
MUX_SEL_UNIT_602 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_557 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_301 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_602
									);
MUX_SEL_UNIT_603 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_813 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_603
									);
MUX_SEL_UNIT_604 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_558 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_302 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_604
									);
MUX_SEL_UNIT_605 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_814 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_605
									);
MUX_SEL_UNIT_606 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_559 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_303 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_606
									);
MUX_SEL_UNIT_607 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_815 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_607
									);
MUX_SEL_UNIT_608 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_560 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_304 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_608
									);
MUX_SEL_UNIT_609 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_816 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_609
									);
MUX_SEL_UNIT_610 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_561 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_305 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_610
									);
MUX_SEL_UNIT_611 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_817 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_611
									);
MUX_SEL_UNIT_612 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_562 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_306 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_612
									);
MUX_SEL_UNIT_613 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_818 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_613
									);
MUX_SEL_UNIT_614 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_563 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_307 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_614
									);
MUX_SEL_UNIT_615 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_819 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_615
									);
MUX_SEL_UNIT_616 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_564 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_308 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_616
									);
MUX_SEL_UNIT_617 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_820 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_617
									);
MUX_SEL_UNIT_618 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_565 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_309 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_618
									);
MUX_SEL_UNIT_619 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_821 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_619
									);
MUX_SEL_UNIT_620 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_566 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_310 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_620
									);
MUX_SEL_UNIT_621 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_822 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_621
									);
MUX_SEL_UNIT_622 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_567 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_311 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_622
									);
MUX_SEL_UNIT_623 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_823 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_623
									);
MUX_SEL_UNIT_624 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_568 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_312 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_624
									);
MUX_SEL_UNIT_625 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_824 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_625
									);
MUX_SEL_UNIT_626 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_569 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_313 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_626
									);
MUX_SEL_UNIT_627 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_825 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_627
									);
MUX_SEL_UNIT_628 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_570 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_314 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_628
									);
MUX_SEL_UNIT_629 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_826 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_629
									);
MUX_SEL_UNIT_630 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_571 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_315 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_630
									);
MUX_SEL_UNIT_631 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_827 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_631
									);
MUX_SEL_UNIT_632 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_572 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_316 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_632
									);
MUX_SEL_UNIT_633 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_828 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_633
									);
MUX_SEL_UNIT_634 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_573 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_317 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_634
									);
MUX_SEL_UNIT_635 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_829 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_635
									);
MUX_SEL_UNIT_636 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_574 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_318 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_636
									);
MUX_SEL_UNIT_637 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_830 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_637
									);
MUX_SEL_UNIT_638 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_575 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_319 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_638
									);
MUX_SEL_UNIT_639 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_831 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_639
									);
MUX_SEL_UNIT_640 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_576 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_320 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_640
									);
MUX_SEL_UNIT_641 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_832 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_641
									);
MUX_SEL_UNIT_642 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_577 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_321 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_642
									);
MUX_SEL_UNIT_643 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_833 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_643
									);
MUX_SEL_UNIT_644 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_578 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_322 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_644
									);
MUX_SEL_UNIT_645 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_834 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_645
									);
MUX_SEL_UNIT_646 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_579 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_323 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_646
									);
MUX_SEL_UNIT_647 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_835 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_647
									);
MUX_SEL_UNIT_648 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_580 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_324 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_648
									);
MUX_SEL_UNIT_649 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_836 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_649
									);
MUX_SEL_UNIT_650 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_581 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_325 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_650
									);
MUX_SEL_UNIT_651 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_837 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_651
									);
MUX_SEL_UNIT_652 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_582 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_326 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_652
									);
MUX_SEL_UNIT_653 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_838 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_653
									);
MUX_SEL_UNIT_654 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_583 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_327 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_654
									);
MUX_SEL_UNIT_655 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_839 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_655
									);
MUX_SEL_UNIT_656 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_584 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_328 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_656
									);
MUX_SEL_UNIT_657 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_840 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_657
									);
MUX_SEL_UNIT_658 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_585 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_329 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_658
									);
MUX_SEL_UNIT_659 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_841 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_659
									);
MUX_SEL_UNIT_660 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_586 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_330 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_660
									);
MUX_SEL_UNIT_661 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_842 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_661
									);
MUX_SEL_UNIT_662 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_587 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_331 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_662
									);
MUX_SEL_UNIT_663 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_843 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_663
									);
MUX_SEL_UNIT_664 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_588 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_332 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_664
									);
MUX_SEL_UNIT_665 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_844 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_665
									);
MUX_SEL_UNIT_666 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_589 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_333 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_666
									);
MUX_SEL_UNIT_667 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_845 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_667
									);
MUX_SEL_UNIT_668 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_590 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_334 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_668
									);
MUX_SEL_UNIT_669 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_846 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_669
									);
MUX_SEL_UNIT_670 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_591 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_335 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_670
									);
MUX_SEL_UNIT_671 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_847 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_671
									);
MUX_SEL_UNIT_672 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_592 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_336 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_672
									);
MUX_SEL_UNIT_673 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_848 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_673
									);
MUX_SEL_UNIT_674 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_593 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_337 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_674
									);
MUX_SEL_UNIT_675 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_849 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_675
									);
MUX_SEL_UNIT_676 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_594 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_338 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_676
									);
MUX_SEL_UNIT_677 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_850 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_677
									);
MUX_SEL_UNIT_678 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_595 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_339 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_678
									);
MUX_SEL_UNIT_679 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_851 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_679
									);
MUX_SEL_UNIT_680 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_596 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_340 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_680
									);
MUX_SEL_UNIT_681 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_852 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_681
									);
MUX_SEL_UNIT_682 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_597 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_341 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_682
									);
MUX_SEL_UNIT_683 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_853 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_683
									);
MUX_SEL_UNIT_684 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_598 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_342 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_684
									);
MUX_SEL_UNIT_685 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_854 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_685
									);
MUX_SEL_UNIT_686 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_599 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_343 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_686
									);
MUX_SEL_UNIT_687 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_855 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_687
									);
MUX_SEL_UNIT_688 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_600 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_344 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_688
									);
MUX_SEL_UNIT_689 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_856 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_689
									);
MUX_SEL_UNIT_690 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_601 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_345 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_690
									);
MUX_SEL_UNIT_691 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_857 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_691
									);
MUX_SEL_UNIT_692 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_602 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_346 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_692
									);
MUX_SEL_UNIT_693 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_858 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_693
									);
MUX_SEL_UNIT_694 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_603 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_347 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_694
									);
MUX_SEL_UNIT_695 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_859 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_695
									);
MUX_SEL_UNIT_696 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_604 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_348 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_696
									);
MUX_SEL_UNIT_697 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_860 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_697
									);
MUX_SEL_UNIT_698 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_605 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_349 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_698
									);
MUX_SEL_UNIT_699 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_861 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_699
									);
MUX_SEL_UNIT_700 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_606 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_350 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_700
									);
MUX_SEL_UNIT_701 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_862 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_701
									);
MUX_SEL_UNIT_702 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_607 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_351 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_702
									);
MUX_SEL_UNIT_703 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_863 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_703
									);
MUX_SEL_UNIT_704 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_608 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_352 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_704
									);
MUX_SEL_UNIT_705 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_864 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_705
									);
MUX_SEL_UNIT_706 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_609 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_353 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_706
									);
MUX_SEL_UNIT_707 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_865 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_707
									);
MUX_SEL_UNIT_708 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_610 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_354 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_708
									);
MUX_SEL_UNIT_709 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_866 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_709
									);
MUX_SEL_UNIT_710 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_611 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_355 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_710
									);
MUX_SEL_UNIT_711 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_867 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_711
									);
MUX_SEL_UNIT_712 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_612 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_356 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_712
									);
MUX_SEL_UNIT_713 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_868 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_713
									);
MUX_SEL_UNIT_714 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_613 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_357 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_714
									);
MUX_SEL_UNIT_715 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_869 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_715
									);
MUX_SEL_UNIT_716 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_614 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_358 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_716
									);
MUX_SEL_UNIT_717 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_870 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_717
									);
MUX_SEL_UNIT_718 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_615 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_359 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_718
									);
MUX_SEL_UNIT_719 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_871 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_719
									);
MUX_SEL_UNIT_720 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_616 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_360 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_720
									);
MUX_SEL_UNIT_721 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_872 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_721
									);
MUX_SEL_UNIT_722 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_617 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_361 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_722
									);
MUX_SEL_UNIT_723 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_873 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_723
									);
MUX_SEL_UNIT_724 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_618 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_362 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_724
									);
MUX_SEL_UNIT_725 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_874 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_725
									);
MUX_SEL_UNIT_726 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_619 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_363 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_726
									);
MUX_SEL_UNIT_727 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_875 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_727
									);
MUX_SEL_UNIT_728 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_620 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_364 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_728
									);
MUX_SEL_UNIT_729 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_876 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_729
									);
MUX_SEL_UNIT_730 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_621 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_365 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_730
									);
MUX_SEL_UNIT_731 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_877 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_731
									);
MUX_SEL_UNIT_732 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_622 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_366 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_732
									);
MUX_SEL_UNIT_733 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_878 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_733
									);
MUX_SEL_UNIT_734 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_623 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_367 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_734
									);
MUX_SEL_UNIT_735 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_879 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_735
									);
MUX_SEL_UNIT_736 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_624 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_368 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_736
									);
MUX_SEL_UNIT_737 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_880 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_737
									);
MUX_SEL_UNIT_738 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_625 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_369 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_738
									);
MUX_SEL_UNIT_739 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_881 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_739
									);
MUX_SEL_UNIT_740 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_626 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_370 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_740
									);
MUX_SEL_UNIT_741 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_882 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_741
									);
MUX_SEL_UNIT_742 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_627 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_371 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_742
									);
MUX_SEL_UNIT_743 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_883 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_743
									);
MUX_SEL_UNIT_744 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_628 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_372 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_744
									);
MUX_SEL_UNIT_745 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_884 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_745
									);
MUX_SEL_UNIT_746 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_629 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_373 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_746
									);
MUX_SEL_UNIT_747 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_885 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_747
									);
MUX_SEL_UNIT_748 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_630 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_374 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_748
									);
MUX_SEL_UNIT_749 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_886 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_749
									);
MUX_SEL_UNIT_750 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_631 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_375 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_750
									);
MUX_SEL_UNIT_751 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_887 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_751
									);
MUX_SEL_UNIT_752 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_632 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_376 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_752
									);
MUX_SEL_UNIT_753 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_888 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_753
									);
MUX_SEL_UNIT_754 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_633 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_377 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_754
									);
MUX_SEL_UNIT_755 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_889 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_755
									);
MUX_SEL_UNIT_756 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_634 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_378 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_756
									);
MUX_SEL_UNIT_757 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_890 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_757
									);
MUX_SEL_UNIT_758 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_635 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_379 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_758
									);
MUX_SEL_UNIT_759 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_891 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_759
									);
MUX_SEL_UNIT_760 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_636 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_380 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_760
									);
MUX_SEL_UNIT_761 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_892 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_761
									);
MUX_SEL_UNIT_762 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_637 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_381 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_762
									);
MUX_SEL_UNIT_763 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_893 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_763
									);
MUX_SEL_UNIT_764 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_638 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_382 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_764
									);
MUX_SEL_UNIT_765 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_894 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_765
									);
MUX_SEL_UNIT_766 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_639 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_383 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_766
									);
MUX_SEL_UNIT_767 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_895 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_767
									);
MUX_SEL_UNIT_768 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_768 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_640 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_384 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_768
									);
MUX_SEL_UNIT_769 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_896 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_769
									);
MUX_SEL_UNIT_770 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_769 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_641 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_385 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_770
									);
MUX_SEL_UNIT_771 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_897 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_771
									);
MUX_SEL_UNIT_772 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_770 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_642 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_386 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_772
									);
MUX_SEL_UNIT_773 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_898 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_773
									);
MUX_SEL_UNIT_774 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_771 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_643 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_387 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_774
									);
MUX_SEL_UNIT_775 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_899 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_775
									);
MUX_SEL_UNIT_776 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_772 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_644 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_388 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_776
									);
MUX_SEL_UNIT_777 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_900 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_777
									);
MUX_SEL_UNIT_778 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_773 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_645 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_389 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_778
									);
MUX_SEL_UNIT_779 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_901 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_779
									);
MUX_SEL_UNIT_780 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_774 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_646 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_390 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_780
									);
MUX_SEL_UNIT_781 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_902 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_781
									);
MUX_SEL_UNIT_782 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_775 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_647 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_391 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_782
									);
MUX_SEL_UNIT_783 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_903 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_783
									);
MUX_SEL_UNIT_784 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_776 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_648 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_392 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_784
									);
MUX_SEL_UNIT_785 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_904 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_785
									);
MUX_SEL_UNIT_786 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_777 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_649 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_393 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_786
									);
MUX_SEL_UNIT_787 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_905 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_787
									);
MUX_SEL_UNIT_788 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_778 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_650 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_394 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_788
									);
MUX_SEL_UNIT_789 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_906 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_789
									);
MUX_SEL_UNIT_790 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_779 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_651 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_395 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_790
									);
MUX_SEL_UNIT_791 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_907 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_791
									);
MUX_SEL_UNIT_792 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_780 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_652 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_396 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_792
									);
MUX_SEL_UNIT_793 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_908 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_793
									);
MUX_SEL_UNIT_794 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_781 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_653 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_397 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_794
									);
MUX_SEL_UNIT_795 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_909 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_795
									);
MUX_SEL_UNIT_796 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_782 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_654 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_398 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_796
									);
MUX_SEL_UNIT_797 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_910 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_797
									);
MUX_SEL_UNIT_798 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_783 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_655 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_399 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_798
									);
MUX_SEL_UNIT_799 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_911 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_799
									);
MUX_SEL_UNIT_800 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_784 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_656 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_400 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_800
									);
MUX_SEL_UNIT_801 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_912 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_801
									);
MUX_SEL_UNIT_802 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_785 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_657 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_401 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_802
									);
MUX_SEL_UNIT_803 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_913 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_803
									);
MUX_SEL_UNIT_804 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_786 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_658 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_402 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_804
									);
MUX_SEL_UNIT_805 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_914 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_805
									);
MUX_SEL_UNIT_806 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_787 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_659 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_403 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_806
									);
MUX_SEL_UNIT_807 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_915 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_807
									);
MUX_SEL_UNIT_808 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_788 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_660 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_404 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_808
									);
MUX_SEL_UNIT_809 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_916 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_809
									);
MUX_SEL_UNIT_810 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_789 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_661 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_405 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_810
									);
MUX_SEL_UNIT_811 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_917 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_811
									);
MUX_SEL_UNIT_812 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_790 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_662 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_406 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_812
									);
MUX_SEL_UNIT_813 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_918 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_813
									);
MUX_SEL_UNIT_814 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_791 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_663 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_407 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_814
									);
MUX_SEL_UNIT_815 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_919 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_815
									);
MUX_SEL_UNIT_816 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_792 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_664 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_408 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_816
									);
MUX_SEL_UNIT_817 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_920 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_817
									);
MUX_SEL_UNIT_818 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_793 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_665 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_409 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_818
									);
MUX_SEL_UNIT_819 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_921 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_819
									);
MUX_SEL_UNIT_820 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_794 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_666 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_410 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_820
									);
MUX_SEL_UNIT_821 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_922 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_821
									);
MUX_SEL_UNIT_822 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_795 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_667 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_411 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_822
									);
MUX_SEL_UNIT_823 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_923 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_823
									);
MUX_SEL_UNIT_824 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_796 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_668 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_412 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_824
									);
MUX_SEL_UNIT_825 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_924 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_825
									);
MUX_SEL_UNIT_826 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_797 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_669 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_413 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_826
									);
MUX_SEL_UNIT_827 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_925 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_827
									);
MUX_SEL_UNIT_828 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_798 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_670 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_414 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_828
									);
MUX_SEL_UNIT_829 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_926 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_829
									);
MUX_SEL_UNIT_830 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_799 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_671 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_415 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_830
									);
MUX_SEL_UNIT_831 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_927 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_831
									);
MUX_SEL_UNIT_832 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_800 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_672 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_416 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_832
									);
MUX_SEL_UNIT_833 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_928 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_833
									);
MUX_SEL_UNIT_834 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_801 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_673 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_417 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_834
									);
MUX_SEL_UNIT_835 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_929 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_835
									);
MUX_SEL_UNIT_836 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_802 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_674 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_418 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_836
									);
MUX_SEL_UNIT_837 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_930 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_837
									);
MUX_SEL_UNIT_838 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_803 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_675 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_419 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_838
									);
MUX_SEL_UNIT_839 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_931 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_839
									);
MUX_SEL_UNIT_840 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_804 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_676 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_420 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_840
									);
MUX_SEL_UNIT_841 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_932 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_841
									);
MUX_SEL_UNIT_842 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_805 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_677 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_421 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_842
									);
MUX_SEL_UNIT_843 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_933 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_843
									);
MUX_SEL_UNIT_844 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_806 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_678 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_422 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_844
									);
MUX_SEL_UNIT_845 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_934 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_845
									);
MUX_SEL_UNIT_846 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_807 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_679 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_423 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_846
									);
MUX_SEL_UNIT_847 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_935 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_847
									);
MUX_SEL_UNIT_848 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_808 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_680 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_424 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_848
									);
MUX_SEL_UNIT_849 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_936 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_849
									);
MUX_SEL_UNIT_850 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_809 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_681 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_425 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_850
									);
MUX_SEL_UNIT_851 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_937 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_851
									);
MUX_SEL_UNIT_852 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_810 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_682 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_426 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_852
									);
MUX_SEL_UNIT_853 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_938 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_853
									);
MUX_SEL_UNIT_854 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_811 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_683 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_427 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_854
									);
MUX_SEL_UNIT_855 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_939 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_855
									);
MUX_SEL_UNIT_856 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_812 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_684 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_428 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_856
									);
MUX_SEL_UNIT_857 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_940 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_857
									);
MUX_SEL_UNIT_858 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_813 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_685 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_429 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_858
									);
MUX_SEL_UNIT_859 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_941 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_859
									);
MUX_SEL_UNIT_860 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_814 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_686 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_430 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_860
									);
MUX_SEL_UNIT_861 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_942 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_861
									);
MUX_SEL_UNIT_862 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_815 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_687 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_431 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_862
									);
MUX_SEL_UNIT_863 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_943 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_863
									);
MUX_SEL_UNIT_864 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_816 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_688 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_432 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_864
									);
MUX_SEL_UNIT_865 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_944 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_865
									);
MUX_SEL_UNIT_866 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_817 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_689 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_433 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_866
									);
MUX_SEL_UNIT_867 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_945 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_867
									);
MUX_SEL_UNIT_868 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_818 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_690 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_434 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_868
									);
MUX_SEL_UNIT_869 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_946 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_869
									);
MUX_SEL_UNIT_870 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_819 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_691 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_435 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_870
									);
MUX_SEL_UNIT_871 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_947 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_871
									);
MUX_SEL_UNIT_872 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_820 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_692 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_436 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_872
									);
MUX_SEL_UNIT_873 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_948 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_873
									);
MUX_SEL_UNIT_874 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_821 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_693 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_437 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_874
									);
MUX_SEL_UNIT_875 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_949 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_875
									);
MUX_SEL_UNIT_876 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_822 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_694 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_438 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_876
									);
MUX_SEL_UNIT_877 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_950 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_877
									);
MUX_SEL_UNIT_878 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_823 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_695 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_439 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_878
									);
MUX_SEL_UNIT_879 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_951 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_879
									);
MUX_SEL_UNIT_880 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_824 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_696 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_440 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_880
									);
MUX_SEL_UNIT_881 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_952 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_881
									);
MUX_SEL_UNIT_882 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_825 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_697 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_441 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_882
									);
MUX_SEL_UNIT_883 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_953 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_883
									);
MUX_SEL_UNIT_884 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_826 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_698 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_442 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_884
									);
MUX_SEL_UNIT_885 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_954 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_885
									);
MUX_SEL_UNIT_886 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_827 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_699 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_443 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_886
									);
MUX_SEL_UNIT_887 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_955 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_887
									);
MUX_SEL_UNIT_888 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_828 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_700 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_444 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_888
									);
MUX_SEL_UNIT_889 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_956 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_889
									);
MUX_SEL_UNIT_890 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_829 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_701 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_445 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_890
									);
MUX_SEL_UNIT_891 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_957 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_891
									);
MUX_SEL_UNIT_892 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_830 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_702 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_446 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_892
									);
MUX_SEL_UNIT_893 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_958 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_893
									);
MUX_SEL_UNIT_894 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_831 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_703 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_447 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_894
									);
MUX_SEL_UNIT_895 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_959 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_895
									);
MUX_SEL_UNIT_896 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_896 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_832 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_704 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_448 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_896
									);
MUX_SEL_UNIT_897 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_960 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_897
									);
MUX_SEL_UNIT_898 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_897 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_833 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_705 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_449 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_898
									);
MUX_SEL_UNIT_899 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_961 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_899
									);
MUX_SEL_UNIT_900 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_898 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_834 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_706 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_450 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_900
									);
MUX_SEL_UNIT_901 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_962 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_901
									);
MUX_SEL_UNIT_902 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_899 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_835 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_707 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_451 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_902
									);
MUX_SEL_UNIT_903 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_963 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_903
									);
MUX_SEL_UNIT_904 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_900 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_836 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_708 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_452 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_904
									);
MUX_SEL_UNIT_905 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_964 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_905
									);
MUX_SEL_UNIT_906 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_901 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_837 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_709 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_453 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_906
									);
MUX_SEL_UNIT_907 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_965 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_907
									);
MUX_SEL_UNIT_908 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_902 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_838 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_710 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_454 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_908
									);
MUX_SEL_UNIT_909 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_966 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_909
									);
MUX_SEL_UNIT_910 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_903 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_839 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_711 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_455 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_910
									);
MUX_SEL_UNIT_911 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_967 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_911
									);
MUX_SEL_UNIT_912 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_904 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_840 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_712 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_456 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_912
									);
MUX_SEL_UNIT_913 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_968 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_913
									);
MUX_SEL_UNIT_914 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_905 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_841 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_713 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_457 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_914
									);
MUX_SEL_UNIT_915 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_969 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_915
									);
MUX_SEL_UNIT_916 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_906 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_842 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_714 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_458 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_916
									);
MUX_SEL_UNIT_917 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_970 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_917
									);
MUX_SEL_UNIT_918 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_907 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_843 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_715 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_459 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_918
									);
MUX_SEL_UNIT_919 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_971 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_919
									);
MUX_SEL_UNIT_920 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_908 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_844 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_716 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_460 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_920
									);
MUX_SEL_UNIT_921 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_972 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_921
									);
MUX_SEL_UNIT_922 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_909 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_845 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_717 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_461 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_922
									);
MUX_SEL_UNIT_923 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_973 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_923
									);
MUX_SEL_UNIT_924 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_910 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_846 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_718 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_462 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_924
									);
MUX_SEL_UNIT_925 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_974 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_925
									);
MUX_SEL_UNIT_926 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_911 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_847 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_719 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_463 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_926
									);
MUX_SEL_UNIT_927 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_975 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_927
									);
MUX_SEL_UNIT_928 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_912 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_848 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_720 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_464 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_928
									);
MUX_SEL_UNIT_929 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_976 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_929
									);
MUX_SEL_UNIT_930 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_913 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_849 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_721 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_465 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_930
									);
MUX_SEL_UNIT_931 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_977 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_931
									);
MUX_SEL_UNIT_932 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_914 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_850 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_722 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_466 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_932
									);
MUX_SEL_UNIT_933 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_978 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_933
									);
MUX_SEL_UNIT_934 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_915 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_851 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_723 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_467 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_934
									);
MUX_SEL_UNIT_935 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_979 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_935
									);
MUX_SEL_UNIT_936 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_916 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_852 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_724 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_468 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_936
									);
MUX_SEL_UNIT_937 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_980 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_937
									);
MUX_SEL_UNIT_938 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_917 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_853 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_725 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_469 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_938
									);
MUX_SEL_UNIT_939 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_981 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_939
									);
MUX_SEL_UNIT_940 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_918 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_854 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_726 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_470 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_940
									);
MUX_SEL_UNIT_941 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_982 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_941
									);
MUX_SEL_UNIT_942 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_919 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_855 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_727 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_471 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_942
									);
MUX_SEL_UNIT_943 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_983 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_943
									);
MUX_SEL_UNIT_944 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_920 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_856 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_728 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_472 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_944
									);
MUX_SEL_UNIT_945 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_984 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_945
									);
MUX_SEL_UNIT_946 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_921 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_857 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_729 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_473 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_946
									);
MUX_SEL_UNIT_947 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_985 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_947
									);
MUX_SEL_UNIT_948 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_922 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_858 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_730 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_474 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_948
									);
MUX_SEL_UNIT_949 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_986 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_949
									);
MUX_SEL_UNIT_950 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_923 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_859 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_731 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_475 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_950
									);
MUX_SEL_UNIT_951 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_987 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_951
									);
MUX_SEL_UNIT_952 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_924 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_860 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_732 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_476 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_952
									);
MUX_SEL_UNIT_953 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_988 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_953
									);
MUX_SEL_UNIT_954 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_925 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_861 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_733 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_477 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_954
									);
MUX_SEL_UNIT_955 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_989 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_955
									);
MUX_SEL_UNIT_956 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_926 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_862 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_734 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_478 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_956
									);
MUX_SEL_UNIT_957 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_990 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_957
									);
MUX_SEL_UNIT_958 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_927 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_863 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_735 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_479 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_958
									);
MUX_SEL_UNIT_959 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_991 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_959
									);
MUX_SEL_UNIT_960 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_960 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_928 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_864 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_736 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_480 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_960
									);
MUX_SEL_UNIT_961 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_992 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_961
									);
MUX_SEL_UNIT_962 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_961 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_929 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_865 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_737 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_481 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_962
									);
MUX_SEL_UNIT_963 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_993 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_963
									);
MUX_SEL_UNIT_964 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_962 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_930 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_866 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_738 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_482 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_964
									);
MUX_SEL_UNIT_965 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_994 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_965
									);
MUX_SEL_UNIT_966 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_963 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_931 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_867 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_739 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_483 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_966
									);
MUX_SEL_UNIT_967 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_995 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_967
									);
MUX_SEL_UNIT_968 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_964 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_932 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_868 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_740 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_484 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_968
									);
MUX_SEL_UNIT_969 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_996 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_969
									);
MUX_SEL_UNIT_970 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_965 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_933 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_869 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_741 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_485 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_970
									);
MUX_SEL_UNIT_971 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_997 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_971
									);
MUX_SEL_UNIT_972 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_966 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_934 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_870 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_742 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_486 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_972
									);
MUX_SEL_UNIT_973 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_998 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_973
									);
MUX_SEL_UNIT_974 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_967 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_935 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_871 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_743 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_487 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_974
									);
MUX_SEL_UNIT_975 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_999 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_975
									);
MUX_SEL_UNIT_976 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_968 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_936 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_872 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_744 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_488 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_976
									);
MUX_SEL_UNIT_977 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1000 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_977
									);
MUX_SEL_UNIT_978 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_969 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_937 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_873 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_745 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_489 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_978
									);
MUX_SEL_UNIT_979 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1001 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_979
									);
MUX_SEL_UNIT_980 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_970 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_938 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_874 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_746 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_490 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_980
									);
MUX_SEL_UNIT_981 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1002 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_981
									);
MUX_SEL_UNIT_982 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_971 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_939 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_875 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_747 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_491 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_982
									);
MUX_SEL_UNIT_983 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1003 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_983
									);
MUX_SEL_UNIT_984 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_972 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_940 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_876 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_748 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_492 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_984
									);
MUX_SEL_UNIT_985 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1004 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_985
									);
MUX_SEL_UNIT_986 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_973 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_941 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_877 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_749 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_493 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_986
									);
MUX_SEL_UNIT_987 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1005 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_987
									);
MUX_SEL_UNIT_988 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_974 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_942 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_878 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_750 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_494 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_988
									);
MUX_SEL_UNIT_989 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1006 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_989
									);
MUX_SEL_UNIT_990 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_975 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_943 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_879 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_751 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_495 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_990
									);
MUX_SEL_UNIT_991 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1007 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_991
									);
MUX_SEL_UNIT_992 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_992 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_976 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_944 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_880 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_752 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_496 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_992
									);
MUX_SEL_UNIT_993 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1008 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_993
									);
MUX_SEL_UNIT_994 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_993 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_977 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_945 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_881 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_753 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_497 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_994
									);
MUX_SEL_UNIT_995 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1009 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_995
									);
MUX_SEL_UNIT_996 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_994 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_978 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_946 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_882 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_754 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_498 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_996
									);
MUX_SEL_UNIT_997 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1010 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_997
									);
MUX_SEL_UNIT_998 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_995 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_979 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_947 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_883 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_755 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_499 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_998
									);
MUX_SEL_UNIT_999 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1011 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_999
									);
MUX_SEL_UNIT_1000 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_996 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_980 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_948 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_884 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_756 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_500 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1000
									);
MUX_SEL_UNIT_1001 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1012 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1001
									);
MUX_SEL_UNIT_1002 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_997 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_981 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_949 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_885 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_757 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_501 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1002
									);
MUX_SEL_UNIT_1003 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1013 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1003
									);
MUX_SEL_UNIT_1004 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_998 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_982 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_950 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_886 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_758 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_502 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1004
									);
MUX_SEL_UNIT_1005 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1014 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1005
									);
MUX_SEL_UNIT_1006 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_999 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_983 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_951 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_887 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_759 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_503 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1006
									);
MUX_SEL_UNIT_1007 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1015 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1007
									);
MUX_SEL_UNIT_1008 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1008 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1000 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_984 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_952 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_888 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_760 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_504 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1008
									);
MUX_SEL_UNIT_1009 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1016 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1009
									);
MUX_SEL_UNIT_1010 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1009 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1001 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_985 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_953 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_889 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_761 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_505 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1010
									);
MUX_SEL_UNIT_1011 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1017 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1011
									);
MUX_SEL_UNIT_1012 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1010 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1002 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_986 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_954 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_890 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_762 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_506 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1012
									);
MUX_SEL_UNIT_1013 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1018 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1013
									);
MUX_SEL_UNIT_1014 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1011 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1003 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_987 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_955 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_891 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_763 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_507 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1014
									);
MUX_SEL_UNIT_1015 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1019 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1015
									);
MUX_SEL_UNIT_1016 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1016 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1012 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1004 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_988 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_956 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_892 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_764 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_508 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1016
									);
MUX_SEL_UNIT_1017 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1020 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1017
									);
MUX_SEL_UNIT_1018 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1017 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1013 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1005 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_989 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_957 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_893 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_765 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_509 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1018
									);
MUX_SEL_UNIT_1019 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1021 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1019
									);
MUX_SEL_UNIT_1020 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1020 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1018 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1014 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1006 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_990 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_958 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_894 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_766 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_510 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1020
									);
MUX_SEL_UNIT_1021 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1022 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1021
									);
MUX_SEL_UNIT_1022 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1022 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1021 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1019 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1015 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1007 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_991 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_959 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_895 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_767 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_511 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1022
									);
MUX_SEL_UNIT_1023 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_1 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_2 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_3 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_4 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_5 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_6 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_7 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_8 => FROM_STATE_REG_1023 ,
										MUX_10_1_IN_9 => FROM_STATE_REG_1023 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => FROM_SELECTION_UNIT_1023
									);

MASKED_INPUT_0 <= FROM_SELECTION_UNIT_0 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_2 <= FROM_SELECTION_UNIT_2 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_4 <= FROM_SELECTION_UNIT_4 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_6 <= FROM_SELECTION_UNIT_6 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_8 <= FROM_SELECTION_UNIT_8 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_10 <= FROM_SELECTION_UNIT_10 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_12 <= FROM_SELECTION_UNIT_12 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_14 <= FROM_SELECTION_UNIT_14 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_16 <= FROM_SELECTION_UNIT_16 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_18 <= FROM_SELECTION_UNIT_18 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_20 <= FROM_SELECTION_UNIT_20 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_22 <= FROM_SELECTION_UNIT_22 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_24 <= FROM_SELECTION_UNIT_24 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_26 <= FROM_SELECTION_UNIT_26 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_28 <= FROM_SELECTION_UNIT_28 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_30 <= FROM_SELECTION_UNIT_30 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_32 <= FROM_SELECTION_UNIT_32 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_34 <= FROM_SELECTION_UNIT_34 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_36 <= FROM_SELECTION_UNIT_36 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_38 <= FROM_SELECTION_UNIT_38 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_40 <= FROM_SELECTION_UNIT_40 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_42 <= FROM_SELECTION_UNIT_42 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_44 <= FROM_SELECTION_UNIT_44 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_46 <= FROM_SELECTION_UNIT_46 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_48 <= FROM_SELECTION_UNIT_48 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_50 <= FROM_SELECTION_UNIT_50 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_52 <= FROM_SELECTION_UNIT_52 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_54 <= FROM_SELECTION_UNIT_54 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_56 <= FROM_SELECTION_UNIT_56 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_58 <= FROM_SELECTION_UNIT_58 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_60 <= FROM_SELECTION_UNIT_60 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_62 <= FROM_SELECTION_UNIT_62 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_64 <= FROM_SELECTION_UNIT_64 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_66 <= FROM_SELECTION_UNIT_66 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_68 <= FROM_SELECTION_UNIT_68 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_70 <= FROM_SELECTION_UNIT_70 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_72 <= FROM_SELECTION_UNIT_72 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_74 <= FROM_SELECTION_UNIT_74 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_76 <= FROM_SELECTION_UNIT_76 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_78 <= FROM_SELECTION_UNIT_78 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_80 <= FROM_SELECTION_UNIT_80 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_82 <= FROM_SELECTION_UNIT_82 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_84 <= FROM_SELECTION_UNIT_84 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_86 <= FROM_SELECTION_UNIT_86 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_88 <= FROM_SELECTION_UNIT_88 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_90 <= FROM_SELECTION_UNIT_90 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_92 <= FROM_SELECTION_UNIT_92 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_94 <= FROM_SELECTION_UNIT_94 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_96 <= FROM_SELECTION_UNIT_96 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_98 <= FROM_SELECTION_UNIT_98 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_100 <= FROM_SELECTION_UNIT_100 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_102 <= FROM_SELECTION_UNIT_102 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_104 <= FROM_SELECTION_UNIT_104 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_106 <= FROM_SELECTION_UNIT_106 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_108 <= FROM_SELECTION_UNIT_108 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_110 <= FROM_SELECTION_UNIT_110 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_112 <= FROM_SELECTION_UNIT_112 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_114 <= FROM_SELECTION_UNIT_114 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_116 <= FROM_SELECTION_UNIT_116 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_118 <= FROM_SELECTION_UNIT_118 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_120 <= FROM_SELECTION_UNIT_120 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_122 <= FROM_SELECTION_UNIT_122 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_124 <= FROM_SELECTION_UNIT_124 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_126 <= FROM_SELECTION_UNIT_126 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_128 <= FROM_SELECTION_UNIT_128 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_130 <= FROM_SELECTION_UNIT_130 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_132 <= FROM_SELECTION_UNIT_132 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_134 <= FROM_SELECTION_UNIT_134 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_136 <= FROM_SELECTION_UNIT_136 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_138 <= FROM_SELECTION_UNIT_138 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_140 <= FROM_SELECTION_UNIT_140 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_142 <= FROM_SELECTION_UNIT_142 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_144 <= FROM_SELECTION_UNIT_144 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_146 <= FROM_SELECTION_UNIT_146 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_148 <= FROM_SELECTION_UNIT_148 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_150 <= FROM_SELECTION_UNIT_150 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_152 <= FROM_SELECTION_UNIT_152 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_154 <= FROM_SELECTION_UNIT_154 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_156 <= FROM_SELECTION_UNIT_156 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_158 <= FROM_SELECTION_UNIT_158 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_160 <= FROM_SELECTION_UNIT_160 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_162 <= FROM_SELECTION_UNIT_162 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_164 <= FROM_SELECTION_UNIT_164 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_166 <= FROM_SELECTION_UNIT_166 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_168 <= FROM_SELECTION_UNIT_168 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_170 <= FROM_SELECTION_UNIT_170 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_172 <= FROM_SELECTION_UNIT_172 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_174 <= FROM_SELECTION_UNIT_174 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_176 <= FROM_SELECTION_UNIT_176 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_178 <= FROM_SELECTION_UNIT_178 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_180 <= FROM_SELECTION_UNIT_180 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_182 <= FROM_SELECTION_UNIT_182 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_184 <= FROM_SELECTION_UNIT_184 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_186 <= FROM_SELECTION_UNIT_186 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_188 <= FROM_SELECTION_UNIT_188 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_190 <= FROM_SELECTION_UNIT_190 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_192 <= FROM_SELECTION_UNIT_192 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_194 <= FROM_SELECTION_UNIT_194 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_196 <= FROM_SELECTION_UNIT_196 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_198 <= FROM_SELECTION_UNIT_198 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_200 <= FROM_SELECTION_UNIT_200 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_202 <= FROM_SELECTION_UNIT_202 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_204 <= FROM_SELECTION_UNIT_204 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_206 <= FROM_SELECTION_UNIT_206 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_208 <= FROM_SELECTION_UNIT_208 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_210 <= FROM_SELECTION_UNIT_210 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_212 <= FROM_SELECTION_UNIT_212 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_214 <= FROM_SELECTION_UNIT_214 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_216 <= FROM_SELECTION_UNIT_216 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_218 <= FROM_SELECTION_UNIT_218 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_220 <= FROM_SELECTION_UNIT_220 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_222 <= FROM_SELECTION_UNIT_222 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_224 <= FROM_SELECTION_UNIT_224 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_226 <= FROM_SELECTION_UNIT_226 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_228 <= FROM_SELECTION_UNIT_228 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_230 <= FROM_SELECTION_UNIT_230 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_232 <= FROM_SELECTION_UNIT_232 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_234 <= FROM_SELECTION_UNIT_234 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_236 <= FROM_SELECTION_UNIT_236 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_238 <= FROM_SELECTION_UNIT_238 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_240 <= FROM_SELECTION_UNIT_240 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_242 <= FROM_SELECTION_UNIT_242 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_244 <= FROM_SELECTION_UNIT_244 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_246 <= FROM_SELECTION_UNIT_246 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_248 <= FROM_SELECTION_UNIT_248 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_250 <= FROM_SELECTION_UNIT_250 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_252 <= FROM_SELECTION_UNIT_252 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_254 <= FROM_SELECTION_UNIT_254 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_256 <= FROM_SELECTION_UNIT_256 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_258 <= FROM_SELECTION_UNIT_258 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_260 <= FROM_SELECTION_UNIT_260 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_262 <= FROM_SELECTION_UNIT_262 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_264 <= FROM_SELECTION_UNIT_264 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_266 <= FROM_SELECTION_UNIT_266 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_268 <= FROM_SELECTION_UNIT_268 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_270 <= FROM_SELECTION_UNIT_270 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_272 <= FROM_SELECTION_UNIT_272 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_274 <= FROM_SELECTION_UNIT_274 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_276 <= FROM_SELECTION_UNIT_276 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_278 <= FROM_SELECTION_UNIT_278 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_280 <= FROM_SELECTION_UNIT_280 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_282 <= FROM_SELECTION_UNIT_282 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_284 <= FROM_SELECTION_UNIT_284 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_286 <= FROM_SELECTION_UNIT_286 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_288 <= FROM_SELECTION_UNIT_288 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_290 <= FROM_SELECTION_UNIT_290 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_292 <= FROM_SELECTION_UNIT_292 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_294 <= FROM_SELECTION_UNIT_294 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_296 <= FROM_SELECTION_UNIT_296 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_298 <= FROM_SELECTION_UNIT_298 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_300 <= FROM_SELECTION_UNIT_300 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_302 <= FROM_SELECTION_UNIT_302 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_304 <= FROM_SELECTION_UNIT_304 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_306 <= FROM_SELECTION_UNIT_306 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_308 <= FROM_SELECTION_UNIT_308 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_310 <= FROM_SELECTION_UNIT_310 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_312 <= FROM_SELECTION_UNIT_312 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_314 <= FROM_SELECTION_UNIT_314 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_316 <= FROM_SELECTION_UNIT_316 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_318 <= FROM_SELECTION_UNIT_318 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_320 <= FROM_SELECTION_UNIT_320 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_322 <= FROM_SELECTION_UNIT_322 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_324 <= FROM_SELECTION_UNIT_324 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_326 <= FROM_SELECTION_UNIT_326 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_328 <= FROM_SELECTION_UNIT_328 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_330 <= FROM_SELECTION_UNIT_330 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_332 <= FROM_SELECTION_UNIT_332 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_334 <= FROM_SELECTION_UNIT_334 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_336 <= FROM_SELECTION_UNIT_336 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_338 <= FROM_SELECTION_UNIT_338 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_340 <= FROM_SELECTION_UNIT_340 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_342 <= FROM_SELECTION_UNIT_342 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_344 <= FROM_SELECTION_UNIT_344 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_346 <= FROM_SELECTION_UNIT_346 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_348 <= FROM_SELECTION_UNIT_348 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_350 <= FROM_SELECTION_UNIT_350 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_352 <= FROM_SELECTION_UNIT_352 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_354 <= FROM_SELECTION_UNIT_354 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_356 <= FROM_SELECTION_UNIT_356 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_358 <= FROM_SELECTION_UNIT_358 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_360 <= FROM_SELECTION_UNIT_360 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_362 <= FROM_SELECTION_UNIT_362 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_364 <= FROM_SELECTION_UNIT_364 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_366 <= FROM_SELECTION_UNIT_366 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_368 <= FROM_SELECTION_UNIT_368 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_370 <= FROM_SELECTION_UNIT_370 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_372 <= FROM_SELECTION_UNIT_372 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_374 <= FROM_SELECTION_UNIT_374 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_376 <= FROM_SELECTION_UNIT_376 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_378 <= FROM_SELECTION_UNIT_378 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_380 <= FROM_SELECTION_UNIT_380 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_382 <= FROM_SELECTION_UNIT_382 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_384 <= FROM_SELECTION_UNIT_384 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_386 <= FROM_SELECTION_UNIT_386 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_388 <= FROM_SELECTION_UNIT_388 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_390 <= FROM_SELECTION_UNIT_390 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_392 <= FROM_SELECTION_UNIT_392 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_394 <= FROM_SELECTION_UNIT_394 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_396 <= FROM_SELECTION_UNIT_396 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_398 <= FROM_SELECTION_UNIT_398 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_400 <= FROM_SELECTION_UNIT_400 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_402 <= FROM_SELECTION_UNIT_402 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_404 <= FROM_SELECTION_UNIT_404 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_406 <= FROM_SELECTION_UNIT_406 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_408 <= FROM_SELECTION_UNIT_408 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_410 <= FROM_SELECTION_UNIT_410 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_412 <= FROM_SELECTION_UNIT_412 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_414 <= FROM_SELECTION_UNIT_414 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_416 <= FROM_SELECTION_UNIT_416 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_418 <= FROM_SELECTION_UNIT_418 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_420 <= FROM_SELECTION_UNIT_420 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_422 <= FROM_SELECTION_UNIT_422 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_424 <= FROM_SELECTION_UNIT_424 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_426 <= FROM_SELECTION_UNIT_426 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_428 <= FROM_SELECTION_UNIT_428 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_430 <= FROM_SELECTION_UNIT_430 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_432 <= FROM_SELECTION_UNIT_432 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_434 <= FROM_SELECTION_UNIT_434 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_436 <= FROM_SELECTION_UNIT_436 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_438 <= FROM_SELECTION_UNIT_438 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_440 <= FROM_SELECTION_UNIT_440 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_442 <= FROM_SELECTION_UNIT_442 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_444 <= FROM_SELECTION_UNIT_444 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_446 <= FROM_SELECTION_UNIT_446 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_448 <= FROM_SELECTION_UNIT_448 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_450 <= FROM_SELECTION_UNIT_450 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_452 <= FROM_SELECTION_UNIT_452 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_454 <= FROM_SELECTION_UNIT_454 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_456 <= FROM_SELECTION_UNIT_456 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_458 <= FROM_SELECTION_UNIT_458 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_460 <= FROM_SELECTION_UNIT_460 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_462 <= FROM_SELECTION_UNIT_462 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_464 <= FROM_SELECTION_UNIT_464 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_466 <= FROM_SELECTION_UNIT_466 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_468 <= FROM_SELECTION_UNIT_468 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_470 <= FROM_SELECTION_UNIT_470 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_472 <= FROM_SELECTION_UNIT_472 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_474 <= FROM_SELECTION_UNIT_474 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_476 <= FROM_SELECTION_UNIT_476 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_478 <= FROM_SELECTION_UNIT_478 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_480 <= FROM_SELECTION_UNIT_480 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_482 <= FROM_SELECTION_UNIT_482 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_484 <= FROM_SELECTION_UNIT_484 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_486 <= FROM_SELECTION_UNIT_486 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_488 <= FROM_SELECTION_UNIT_488 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_490 <= FROM_SELECTION_UNIT_490 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_492 <= FROM_SELECTION_UNIT_492 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_494 <= FROM_SELECTION_UNIT_494 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_496 <= FROM_SELECTION_UNIT_496 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_498 <= FROM_SELECTION_UNIT_498 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_500 <= FROM_SELECTION_UNIT_500 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_502 <= FROM_SELECTION_UNIT_502 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_504 <= FROM_SELECTION_UNIT_504 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_506 <= FROM_SELECTION_UNIT_506 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_508 <= FROM_SELECTION_UNIT_508 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_510 <= FROM_SELECTION_UNIT_510 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_512 <= FROM_SELECTION_UNIT_512 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_514 <= FROM_SELECTION_UNIT_514 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_516 <= FROM_SELECTION_UNIT_516 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_518 <= FROM_SELECTION_UNIT_518 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_520 <= FROM_SELECTION_UNIT_520 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_522 <= FROM_SELECTION_UNIT_522 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_524 <= FROM_SELECTION_UNIT_524 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_526 <= FROM_SELECTION_UNIT_526 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_528 <= FROM_SELECTION_UNIT_528 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_530 <= FROM_SELECTION_UNIT_530 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_532 <= FROM_SELECTION_UNIT_532 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_534 <= FROM_SELECTION_UNIT_534 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_536 <= FROM_SELECTION_UNIT_536 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_538 <= FROM_SELECTION_UNIT_538 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_540 <= FROM_SELECTION_UNIT_540 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_542 <= FROM_SELECTION_UNIT_542 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_544 <= FROM_SELECTION_UNIT_544 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_546 <= FROM_SELECTION_UNIT_546 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_548 <= FROM_SELECTION_UNIT_548 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_550 <= FROM_SELECTION_UNIT_550 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_552 <= FROM_SELECTION_UNIT_552 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_554 <= FROM_SELECTION_UNIT_554 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_556 <= FROM_SELECTION_UNIT_556 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_558 <= FROM_SELECTION_UNIT_558 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_560 <= FROM_SELECTION_UNIT_560 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_562 <= FROM_SELECTION_UNIT_562 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_564 <= FROM_SELECTION_UNIT_564 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_566 <= FROM_SELECTION_UNIT_566 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_568 <= FROM_SELECTION_UNIT_568 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_570 <= FROM_SELECTION_UNIT_570 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_572 <= FROM_SELECTION_UNIT_572 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_574 <= FROM_SELECTION_UNIT_574 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_576 <= FROM_SELECTION_UNIT_576 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_578 <= FROM_SELECTION_UNIT_578 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_580 <= FROM_SELECTION_UNIT_580 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_582 <= FROM_SELECTION_UNIT_582 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_584 <= FROM_SELECTION_UNIT_584 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_586 <= FROM_SELECTION_UNIT_586 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_588 <= FROM_SELECTION_UNIT_588 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_590 <= FROM_SELECTION_UNIT_590 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_592 <= FROM_SELECTION_UNIT_592 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_594 <= FROM_SELECTION_UNIT_594 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_596 <= FROM_SELECTION_UNIT_596 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_598 <= FROM_SELECTION_UNIT_598 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_600 <= FROM_SELECTION_UNIT_600 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_602 <= FROM_SELECTION_UNIT_602 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_604 <= FROM_SELECTION_UNIT_604 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_606 <= FROM_SELECTION_UNIT_606 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_608 <= FROM_SELECTION_UNIT_608 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_610 <= FROM_SELECTION_UNIT_610 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_612 <= FROM_SELECTION_UNIT_612 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_614 <= FROM_SELECTION_UNIT_614 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_616 <= FROM_SELECTION_UNIT_616 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_618 <= FROM_SELECTION_UNIT_618 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_620 <= FROM_SELECTION_UNIT_620 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_622 <= FROM_SELECTION_UNIT_622 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_624 <= FROM_SELECTION_UNIT_624 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_626 <= FROM_SELECTION_UNIT_626 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_628 <= FROM_SELECTION_UNIT_628 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_630 <= FROM_SELECTION_UNIT_630 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_632 <= FROM_SELECTION_UNIT_632 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_634 <= FROM_SELECTION_UNIT_634 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_636 <= FROM_SELECTION_UNIT_636 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_638 <= FROM_SELECTION_UNIT_638 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_640 <= FROM_SELECTION_UNIT_640 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_642 <= FROM_SELECTION_UNIT_642 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_644 <= FROM_SELECTION_UNIT_644 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_646 <= FROM_SELECTION_UNIT_646 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_648 <= FROM_SELECTION_UNIT_648 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_650 <= FROM_SELECTION_UNIT_650 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_652 <= FROM_SELECTION_UNIT_652 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_654 <= FROM_SELECTION_UNIT_654 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_656 <= FROM_SELECTION_UNIT_656 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_658 <= FROM_SELECTION_UNIT_658 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_660 <= FROM_SELECTION_UNIT_660 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_662 <= FROM_SELECTION_UNIT_662 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_664 <= FROM_SELECTION_UNIT_664 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_666 <= FROM_SELECTION_UNIT_666 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_668 <= FROM_SELECTION_UNIT_668 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_670 <= FROM_SELECTION_UNIT_670 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_672 <= FROM_SELECTION_UNIT_672 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_674 <= FROM_SELECTION_UNIT_674 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_676 <= FROM_SELECTION_UNIT_676 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_678 <= FROM_SELECTION_UNIT_678 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_680 <= FROM_SELECTION_UNIT_680 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_682 <= FROM_SELECTION_UNIT_682 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_684 <= FROM_SELECTION_UNIT_684 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_686 <= FROM_SELECTION_UNIT_686 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_688 <= FROM_SELECTION_UNIT_688 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_690 <= FROM_SELECTION_UNIT_690 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_692 <= FROM_SELECTION_UNIT_692 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_694 <= FROM_SELECTION_UNIT_694 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_696 <= FROM_SELECTION_UNIT_696 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_698 <= FROM_SELECTION_UNIT_698 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_700 <= FROM_SELECTION_UNIT_700 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_702 <= FROM_SELECTION_UNIT_702 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_704 <= FROM_SELECTION_UNIT_704 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_706 <= FROM_SELECTION_UNIT_706 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_708 <= FROM_SELECTION_UNIT_708 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_710 <= FROM_SELECTION_UNIT_710 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_712 <= FROM_SELECTION_UNIT_712 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_714 <= FROM_SELECTION_UNIT_714 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_716 <= FROM_SELECTION_UNIT_716 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_718 <= FROM_SELECTION_UNIT_718 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_720 <= FROM_SELECTION_UNIT_720 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_722 <= FROM_SELECTION_UNIT_722 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_724 <= FROM_SELECTION_UNIT_724 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_726 <= FROM_SELECTION_UNIT_726 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_728 <= FROM_SELECTION_UNIT_728 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_730 <= FROM_SELECTION_UNIT_730 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_732 <= FROM_SELECTION_UNIT_732 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_734 <= FROM_SELECTION_UNIT_734 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_736 <= FROM_SELECTION_UNIT_736 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_738 <= FROM_SELECTION_UNIT_738 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_740 <= FROM_SELECTION_UNIT_740 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_742 <= FROM_SELECTION_UNIT_742 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_744 <= FROM_SELECTION_UNIT_744 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_746 <= FROM_SELECTION_UNIT_746 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_748 <= FROM_SELECTION_UNIT_748 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_750 <= FROM_SELECTION_UNIT_750 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_752 <= FROM_SELECTION_UNIT_752 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_754 <= FROM_SELECTION_UNIT_754 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_756 <= FROM_SELECTION_UNIT_756 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_758 <= FROM_SELECTION_UNIT_758 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_760 <= FROM_SELECTION_UNIT_760 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_762 <= FROM_SELECTION_UNIT_762 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_764 <= FROM_SELECTION_UNIT_764 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_766 <= FROM_SELECTION_UNIT_766 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_768 <= FROM_SELECTION_UNIT_768 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_770 <= FROM_SELECTION_UNIT_770 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_772 <= FROM_SELECTION_UNIT_772 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_774 <= FROM_SELECTION_UNIT_774 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_776 <= FROM_SELECTION_UNIT_776 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_778 <= FROM_SELECTION_UNIT_778 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_780 <= FROM_SELECTION_UNIT_780 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_782 <= FROM_SELECTION_UNIT_782 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_784 <= FROM_SELECTION_UNIT_784 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_786 <= FROM_SELECTION_UNIT_786 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_788 <= FROM_SELECTION_UNIT_788 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_790 <= FROM_SELECTION_UNIT_790 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_792 <= FROM_SELECTION_UNIT_792 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_794 <= FROM_SELECTION_UNIT_794 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_796 <= FROM_SELECTION_UNIT_796 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_798 <= FROM_SELECTION_UNIT_798 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_800 <= FROM_SELECTION_UNIT_800 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_802 <= FROM_SELECTION_UNIT_802 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_804 <= FROM_SELECTION_UNIT_804 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_806 <= FROM_SELECTION_UNIT_806 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_808 <= FROM_SELECTION_UNIT_808 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_810 <= FROM_SELECTION_UNIT_810 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_812 <= FROM_SELECTION_UNIT_812 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_814 <= FROM_SELECTION_UNIT_814 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_816 <= FROM_SELECTION_UNIT_816 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_818 <= FROM_SELECTION_UNIT_818 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_820 <= FROM_SELECTION_UNIT_820 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_822 <= FROM_SELECTION_UNIT_822 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_824 <= FROM_SELECTION_UNIT_824 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_826 <= FROM_SELECTION_UNIT_826 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_828 <= FROM_SELECTION_UNIT_828 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_830 <= FROM_SELECTION_UNIT_830 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_832 <= FROM_SELECTION_UNIT_832 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_834 <= FROM_SELECTION_UNIT_834 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_836 <= FROM_SELECTION_UNIT_836 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_838 <= FROM_SELECTION_UNIT_838 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_840 <= FROM_SELECTION_UNIT_840 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_842 <= FROM_SELECTION_UNIT_842 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_844 <= FROM_SELECTION_UNIT_844 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_846 <= FROM_SELECTION_UNIT_846 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_848 <= FROM_SELECTION_UNIT_848 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_850 <= FROM_SELECTION_UNIT_850 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_852 <= FROM_SELECTION_UNIT_852 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_854 <= FROM_SELECTION_UNIT_854 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_856 <= FROM_SELECTION_UNIT_856 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_858 <= FROM_SELECTION_UNIT_858 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_860 <= FROM_SELECTION_UNIT_860 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_862 <= FROM_SELECTION_UNIT_862 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_864 <= FROM_SELECTION_UNIT_864 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_866 <= FROM_SELECTION_UNIT_866 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_868 <= FROM_SELECTION_UNIT_868 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_870 <= FROM_SELECTION_UNIT_870 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_872 <= FROM_SELECTION_UNIT_872 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_874 <= FROM_SELECTION_UNIT_874 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_876 <= FROM_SELECTION_UNIT_876 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_878 <= FROM_SELECTION_UNIT_878 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_880 <= FROM_SELECTION_UNIT_880 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_882 <= FROM_SELECTION_UNIT_882 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_884 <= FROM_SELECTION_UNIT_884 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_886 <= FROM_SELECTION_UNIT_886 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_888 <= FROM_SELECTION_UNIT_888 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_890 <= FROM_SELECTION_UNIT_890 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_892 <= FROM_SELECTION_UNIT_892 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_894 <= FROM_SELECTION_UNIT_894 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_896 <= FROM_SELECTION_UNIT_896 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_898 <= FROM_SELECTION_UNIT_898 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_900 <= FROM_SELECTION_UNIT_900 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_902 <= FROM_SELECTION_UNIT_902 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_904 <= FROM_SELECTION_UNIT_904 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_906 <= FROM_SELECTION_UNIT_906 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_908 <= FROM_SELECTION_UNIT_908 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_910 <= FROM_SELECTION_UNIT_910 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_912 <= FROM_SELECTION_UNIT_912 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_914 <= FROM_SELECTION_UNIT_914 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_916 <= FROM_SELECTION_UNIT_916 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_918 <= FROM_SELECTION_UNIT_918 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_920 <= FROM_SELECTION_UNIT_920 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_922 <= FROM_SELECTION_UNIT_922 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_924 <= FROM_SELECTION_UNIT_924 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_926 <= FROM_SELECTION_UNIT_926 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_928 <= FROM_SELECTION_UNIT_928 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_930 <= FROM_SELECTION_UNIT_930 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_932 <= FROM_SELECTION_UNIT_932 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_934 <= FROM_SELECTION_UNIT_934 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_936 <= FROM_SELECTION_UNIT_936 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_938 <= FROM_SELECTION_UNIT_938 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_940 <= FROM_SELECTION_UNIT_940 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_942 <= FROM_SELECTION_UNIT_942 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_944 <= FROM_SELECTION_UNIT_944 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_946 <= FROM_SELECTION_UNIT_946 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_948 <= FROM_SELECTION_UNIT_948 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_950 <= FROM_SELECTION_UNIT_950 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_952 <= FROM_SELECTION_UNIT_952 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_954 <= FROM_SELECTION_UNIT_954 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_956 <= FROM_SELECTION_UNIT_956 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_958 <= FROM_SELECTION_UNIT_958 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_960 <= FROM_SELECTION_UNIT_960 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_962 <= FROM_SELECTION_UNIT_962 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_964 <= FROM_SELECTION_UNIT_964 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_966 <= FROM_SELECTION_UNIT_966 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_968 <= FROM_SELECTION_UNIT_968 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_970 <= FROM_SELECTION_UNIT_970 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_972 <= FROM_SELECTION_UNIT_972 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_974 <= FROM_SELECTION_UNIT_974 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_976 <= FROM_SELECTION_UNIT_976 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_978 <= FROM_SELECTION_UNIT_978 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_980 <= FROM_SELECTION_UNIT_980 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_982 <= FROM_SELECTION_UNIT_982 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_984 <= FROM_SELECTION_UNIT_984 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_986 <= FROM_SELECTION_UNIT_986 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_988 <= FROM_SELECTION_UNIT_988 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_990 <= FROM_SELECTION_UNIT_990 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_992 <= FROM_SELECTION_UNIT_992 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_994 <= FROM_SELECTION_UNIT_994 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_996 <= FROM_SELECTION_UNIT_996 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_998 <= FROM_SELECTION_UNIT_998 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1000 <= FROM_SELECTION_UNIT_1000 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1002 <= FROM_SELECTION_UNIT_1002 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1004 <= FROM_SELECTION_UNIT_1004 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1006 <= FROM_SELECTION_UNIT_1006 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1008 <= FROM_SELECTION_UNIT_1008 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1010 <= FROM_SELECTION_UNIT_1010 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1012 <= FROM_SELECTION_UNIT_1012 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1014 <= FROM_SELECTION_UNIT_1014 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1016 <= FROM_SELECTION_UNIT_1016 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1018 <= FROM_SELECTION_UNIT_1018 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1020 <= FROM_SELECTION_UNIT_1020 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_1022 <= FROM_SELECTION_UNIT_1022 WHEN QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');

FROM_WINDOW_DEC_MASK <= "1";

UNWINDOWED_MASK(0) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(2) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(3) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(4) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(5) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(6) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(7) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(8) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(9) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(10) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(11) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(12) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(13) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(14) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(15) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(16) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(17) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(18) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(19) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(20) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(21) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(22) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(23) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(24) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(25) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(26) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(27) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(28) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(29) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(30) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(31) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(32) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(33) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(34) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(35) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(36) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(37) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(38) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(39) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(40) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(41) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(42) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(43) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(44) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(45) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(46) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(47) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(48) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(49) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(50) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(51) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(52) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(53) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(54) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(55) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(56) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(57) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(58) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(59) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(60) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(61) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(62) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(63) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(64) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(65) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(66) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(67) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(68) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(69) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(70) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(71) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(72) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(73) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(74) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(75) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(76) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(77) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(78) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(79) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(80) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(81) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(82) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(83) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(84) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(85) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(86) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(87) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(88) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(89) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(90) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(91) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(92) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(93) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(94) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(95) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(96) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(97) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(98) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(99) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(100) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(101) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(102) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(103) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(104) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(105) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(106) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(107) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(108) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(109) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(110) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(111) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(112) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(113) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(114) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(115) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(116) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(117) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(118) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(119) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(120) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(121) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(122) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(123) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(124) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(125) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(126) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(127) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(128) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(129) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(130) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(131) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(132) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(133) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(134) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(135) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(136) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(137) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(138) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(139) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(140) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(141) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(142) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(143) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(144) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(145) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(146) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(147) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(148) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(149) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(150) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(151) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(152) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(153) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(154) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(155) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(156) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(157) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(158) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(159) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(160) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(161) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(162) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(163) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(164) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(165) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(166) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(167) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(168) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(169) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(170) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(171) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(172) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(173) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(174) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(175) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(176) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(177) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(178) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(179) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(180) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(181) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(182) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(183) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(184) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(185) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(186) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(187) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(188) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(189) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(190) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(191) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(192) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(193) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(194) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(195) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(196) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(197) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(198) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(199) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(200) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(201) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(202) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(203) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(204) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(205) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(206) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(207) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(208) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(209) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(210) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(211) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(212) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(213) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(214) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(215) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(216) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(217) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(218) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(219) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(220) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(221) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(222) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(223) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(224) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(225) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(226) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(227) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(228) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(229) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(230) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(231) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(232) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(233) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(234) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(235) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(236) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(237) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(238) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(239) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(240) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(241) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(242) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(243) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(244) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(245) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(246) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(247) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(248) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(249) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(250) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(251) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(252) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(253) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(254) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(255) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(256) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(257) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(258) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(259) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(260) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(261) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(262) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(263) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(264) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(265) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(266) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(267) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(268) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(269) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(270) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(271) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(272) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(273) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(274) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(275) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(276) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(277) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(278) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(279) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(280) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(281) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(282) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(283) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(284) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(285) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(286) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(287) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(288) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(289) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(290) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(291) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(292) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(293) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(294) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(295) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(296) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(297) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(298) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(299) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(300) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(301) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(302) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(303) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(304) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(305) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(306) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(307) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(308) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(309) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(310) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(311) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(312) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(313) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(314) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(315) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(316) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(317) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(318) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(319) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(320) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(321) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(322) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(323) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(324) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(325) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(326) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(327) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(328) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(329) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(330) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(331) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(332) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(333) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(334) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(335) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(336) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(337) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(338) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(339) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(340) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(341) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(342) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(343) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(344) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(345) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(346) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(347) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(348) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(349) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(350) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(351) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(352) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(353) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(354) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(355) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(356) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(357) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(358) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(359) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(360) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(361) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(362) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(363) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(364) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(365) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(366) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(367) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(368) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(369) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(370) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(371) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(372) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(373) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(374) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(375) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(376) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(377) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(378) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(379) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(380) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(381) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(382) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(383) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(384) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(385) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(386) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(387) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(388) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(389) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(390) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(391) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(392) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(393) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(394) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(395) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(396) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(397) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(398) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(399) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(400) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(401) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(402) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(403) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(404) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(405) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(406) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(407) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(408) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(409) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(410) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(411) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(412) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(413) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(414) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(415) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(416) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(417) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(418) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(419) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(420) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(421) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(422) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(423) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(424) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(425) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(426) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(427) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(428) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(429) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(430) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(431) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(432) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(433) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(434) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(435) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(436) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(437) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(438) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(439) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(440) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(441) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(442) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(443) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(444) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(445) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(446) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(447) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(448) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(449) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(450) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(451) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(452) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(453) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(454) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(455) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(456) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(457) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(458) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(459) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(460) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(461) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(462) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(463) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(464) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(465) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(466) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(467) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(468) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(469) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(470) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(471) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(472) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(473) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(474) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(475) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(476) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(477) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(478) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(479) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(480) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(481) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(482) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(483) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(484) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(485) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(486) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(487) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(488) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(489) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(490) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(491) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(492) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(493) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(494) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(495) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(496) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(497) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(498) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(499) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(500) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(501) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(502) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(503) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(504) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(505) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(506) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(507) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(508) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(509) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(510) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(511) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(512) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(513) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(514) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(515) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(516) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(517) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(518) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(519) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(520) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(521) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(522) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(523) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(524) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(525) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(526) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(527) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(528) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(529) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(530) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(531) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(532) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(533) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(534) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(535) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(536) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(537) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(538) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(539) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(540) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(541) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(542) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(543) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(544) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(545) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(546) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(547) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(548) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(549) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(550) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(551) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(552) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(553) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(554) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(555) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(556) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(557) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(558) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(559) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(560) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(561) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(562) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(563) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(564) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(565) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(566) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(567) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(568) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(569) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(570) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(571) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(572) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(573) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(574) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(575) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(576) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(577) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(578) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(579) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(580) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(581) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(582) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(583) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(584) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(585) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(586) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(587) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(588) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(589) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(590) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(591) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(592) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(593) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(594) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(595) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(596) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(597) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(598) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(599) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(600) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(601) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(602) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(603) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(604) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(605) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(606) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(607) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(608) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(609) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(610) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(611) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(612) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(613) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(614) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(615) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(616) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(617) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(618) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(619) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(620) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(621) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(622) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(623) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(624) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(625) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(626) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(627) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(628) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(629) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(630) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(631) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(632) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(633) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(634) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(635) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(636) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(637) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(638) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(639) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(640) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(641) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(642) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(643) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(644) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(645) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(646) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(647) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(648) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(649) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(650) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(651) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(652) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(653) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(654) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(655) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(656) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(657) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(658) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(659) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(660) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(661) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(662) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(663) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(664) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(665) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(666) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(667) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(668) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(669) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(670) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(671) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(672) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(673) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(674) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(675) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(676) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(677) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(678) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(679) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(680) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(681) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(682) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(683) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(684) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(685) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(686) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(687) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(688) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(689) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(690) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(691) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(692) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(693) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(694) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(695) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(696) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(697) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(698) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(699) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(700) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(701) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(702) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(703) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(704) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(705) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(706) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(707) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(708) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(709) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(710) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(711) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(712) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(713) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(714) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(715) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(716) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(717) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(718) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(719) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(720) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(721) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(722) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(723) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(724) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(725) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(726) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(727) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(728) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(729) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(730) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(731) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(732) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(733) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(734) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(735) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(736) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(737) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(738) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(739) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(740) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(741) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(742) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(743) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(744) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(745) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(746) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(747) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(748) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(749) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(750) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(751) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(752) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(753) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(754) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(755) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(756) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(757) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(758) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(759) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(760) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(761) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(762) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(763) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(764) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(765) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(766) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(767) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(768) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(769) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(770) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(771) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(772) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(773) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(774) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(775) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(776) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(777) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(778) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(779) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(780) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(781) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(782) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(783) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(784) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(785) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(786) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(787) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(788) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(789) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(790) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(791) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(792) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(793) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(794) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(795) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(796) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(797) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(798) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(799) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(800) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(801) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(802) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(803) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(804) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(805) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(806) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(807) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(808) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(809) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(810) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(811) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(812) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(813) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(814) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(815) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(816) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(817) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(818) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(819) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(820) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(821) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(822) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(823) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(824) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(825) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(826) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(827) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(828) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(829) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(830) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(831) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(832) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(833) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(834) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(835) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(836) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(837) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(838) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(839) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(840) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(841) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(842) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(843) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(844) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(845) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(846) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(847) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(848) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(849) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(850) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(851) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(852) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(853) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(854) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(855) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(856) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(857) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(858) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(859) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(860) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(861) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(862) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(863) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(864) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(865) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(866) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(867) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(868) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(869) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(870) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(871) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(872) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(873) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(874) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(875) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(876) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(877) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(878) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(879) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(880) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(881) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(882) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(883) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(884) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(885) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(886) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(887) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(888) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(889) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(890) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(891) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(892) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(893) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(894) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(895) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(896) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(897) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(898) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(899) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(900) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(901) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(902) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(903) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(904) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(905) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(906) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(907) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(908) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(909) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(910) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(911) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(912) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(913) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(914) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(915) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(916) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(917) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(918) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(919) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(920) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(921) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(922) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(923) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(924) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(925) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(926) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(927) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(928) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(929) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(930) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(931) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(932) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(933) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(934) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(935) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(936) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(937) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(938) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(939) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(940) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(941) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(942) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(943) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(944) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(945) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(946) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(947) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(948) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(949) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(950) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(951) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(952) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(953) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(954) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(955) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(956) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(957) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(958) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(959) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(960) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(961) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(962) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(963) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(964) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(965) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(966) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(967) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(968) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(969) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(970) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(971) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(972) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(973) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(974) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(975) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(976) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(977) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(978) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(979) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(980) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(981) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(982) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(983) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(984) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(985) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(986) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(987) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(988) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(989) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(990) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(991) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(992) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(993) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(994) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(995) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(996) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(997) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(998) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(999) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1000) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1001) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1002) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1003) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1004) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1005) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1006) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1007) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1008) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1009) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1010) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1011) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1012) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1013) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1014) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1015) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1016) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1017) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1018) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1019) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1020) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1021) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1022) <= QEP_N_10_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1023) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1023) <= FROM_WINDOW_DEC_MASK(0);
MUX_REORD_UPDATE_0 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(0 DOWNTO 0) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(0 DOWNTO 0)
									);
MUX_REORD_UPDATE_1 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(2 DOWNTO 2) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1 DOWNTO 1)
									);
MUX_REORD_UPDATE_2 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(4 DOWNTO 4) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(2 DOWNTO 2)
									);
MUX_REORD_UPDATE_3 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(6 DOWNTO 6) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(3 DOWNTO 3)
									);
MUX_REORD_UPDATE_4 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(8 DOWNTO 8) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(4 DOWNTO 4)
									);
MUX_REORD_UPDATE_5 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(10 DOWNTO 10) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(5 DOWNTO 5)
									);
MUX_REORD_UPDATE_6 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(12 DOWNTO 12) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(6 DOWNTO 6)
									);
MUX_REORD_UPDATE_7 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(14 DOWNTO 14) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(7 DOWNTO 7)
									);
MUX_REORD_UPDATE_8 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(16 DOWNTO 16) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(8 DOWNTO 8)
									);
MUX_REORD_UPDATE_9 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(18 DOWNTO 18) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(9 DOWNTO 9)
									);
MUX_REORD_UPDATE_10 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(20 DOWNTO 20) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(10 DOWNTO 10)
									);
MUX_REORD_UPDATE_11 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(22 DOWNTO 22) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(11 DOWNTO 11)
									);
MUX_REORD_UPDATE_12 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(24 DOWNTO 24) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(12 DOWNTO 12)
									);
MUX_REORD_UPDATE_13 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(26 DOWNTO 26) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(13 DOWNTO 13)
									);
MUX_REORD_UPDATE_14 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(28 DOWNTO 28) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(14 DOWNTO 14)
									);
MUX_REORD_UPDATE_15 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(30 DOWNTO 30) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(15 DOWNTO 15)
									);
MUX_REORD_UPDATE_16 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(32 DOWNTO 32) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(16 DOWNTO 16)
									);
MUX_REORD_UPDATE_17 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(34 DOWNTO 34) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(17 DOWNTO 17)
									);
MUX_REORD_UPDATE_18 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(36 DOWNTO 36) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(18 DOWNTO 18)
									);
MUX_REORD_UPDATE_19 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(38 DOWNTO 38) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(19 DOWNTO 19)
									);
MUX_REORD_UPDATE_20 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(40 DOWNTO 40) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(20 DOWNTO 20)
									);
MUX_REORD_UPDATE_21 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(42 DOWNTO 42) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(21 DOWNTO 21)
									);
MUX_REORD_UPDATE_22 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(44 DOWNTO 44) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(22 DOWNTO 22)
									);
MUX_REORD_UPDATE_23 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(46 DOWNTO 46) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(23 DOWNTO 23)
									);
MUX_REORD_UPDATE_24 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(48 DOWNTO 48) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(24 DOWNTO 24)
									);
MUX_REORD_UPDATE_25 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(50 DOWNTO 50) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(25 DOWNTO 25)
									);
MUX_REORD_UPDATE_26 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(52 DOWNTO 52) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(26 DOWNTO 26)
									);
MUX_REORD_UPDATE_27 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(54 DOWNTO 54) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(27 DOWNTO 27)
									);
MUX_REORD_UPDATE_28 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(56 DOWNTO 56) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(28 DOWNTO 28)
									);
MUX_REORD_UPDATE_29 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(58 DOWNTO 58) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(29 DOWNTO 29)
									);
MUX_REORD_UPDATE_30 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(60 DOWNTO 60) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(30 DOWNTO 30)
									);
MUX_REORD_UPDATE_31 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(62 DOWNTO 62) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(31 DOWNTO 31)
									);
MUX_REORD_UPDATE_32 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(64 DOWNTO 64) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(32 DOWNTO 32)
									);
MUX_REORD_UPDATE_33 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(66 DOWNTO 66) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(33 DOWNTO 33)
									);
MUX_REORD_UPDATE_34 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(68 DOWNTO 68) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(34 DOWNTO 34)
									);
MUX_REORD_UPDATE_35 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(70 DOWNTO 70) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(35 DOWNTO 35)
									);
MUX_REORD_UPDATE_36 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(72 DOWNTO 72) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(36 DOWNTO 36)
									);
MUX_REORD_UPDATE_37 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(74 DOWNTO 74) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(37 DOWNTO 37)
									);
MUX_REORD_UPDATE_38 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(76 DOWNTO 76) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(38 DOWNTO 38)
									);
MUX_REORD_UPDATE_39 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(78 DOWNTO 78) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(39 DOWNTO 39)
									);
MUX_REORD_UPDATE_40 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(80 DOWNTO 80) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(40 DOWNTO 40)
									);
MUX_REORD_UPDATE_41 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(82 DOWNTO 82) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(41 DOWNTO 41)
									);
MUX_REORD_UPDATE_42 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(84 DOWNTO 84) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(42 DOWNTO 42)
									);
MUX_REORD_UPDATE_43 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(86 DOWNTO 86) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(43 DOWNTO 43)
									);
MUX_REORD_UPDATE_44 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(88 DOWNTO 88) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(44 DOWNTO 44)
									);
MUX_REORD_UPDATE_45 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(90 DOWNTO 90) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(45 DOWNTO 45)
									);
MUX_REORD_UPDATE_46 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(92 DOWNTO 92) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(46 DOWNTO 46)
									);
MUX_REORD_UPDATE_47 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(94 DOWNTO 94) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(47 DOWNTO 47)
									);
MUX_REORD_UPDATE_48 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(96 DOWNTO 96) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(48 DOWNTO 48)
									);
MUX_REORD_UPDATE_49 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(98 DOWNTO 98) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(49 DOWNTO 49)
									);
MUX_REORD_UPDATE_50 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(100 DOWNTO 100) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(50 DOWNTO 50)
									);
MUX_REORD_UPDATE_51 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(102 DOWNTO 102) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(51 DOWNTO 51)
									);
MUX_REORD_UPDATE_52 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(104 DOWNTO 104) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(52 DOWNTO 52)
									);
MUX_REORD_UPDATE_53 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(106 DOWNTO 106) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(53 DOWNTO 53)
									);
MUX_REORD_UPDATE_54 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(108 DOWNTO 108) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(54 DOWNTO 54)
									);
MUX_REORD_UPDATE_55 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(110 DOWNTO 110) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(55 DOWNTO 55)
									);
MUX_REORD_UPDATE_56 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(112 DOWNTO 112) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(56 DOWNTO 56)
									);
MUX_REORD_UPDATE_57 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(114 DOWNTO 114) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(57 DOWNTO 57)
									);
MUX_REORD_UPDATE_58 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(116 DOWNTO 116) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(58 DOWNTO 58)
									);
MUX_REORD_UPDATE_59 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(118 DOWNTO 118) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(59 DOWNTO 59)
									);
MUX_REORD_UPDATE_60 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(120 DOWNTO 120) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(60 DOWNTO 60)
									);
MUX_REORD_UPDATE_61 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(122 DOWNTO 122) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(61 DOWNTO 61)
									);
MUX_REORD_UPDATE_62 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(124 DOWNTO 124) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(62 DOWNTO 62)
									);
MUX_REORD_UPDATE_63 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(126 DOWNTO 126) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(63 DOWNTO 63)
									);
MUX_REORD_UPDATE_64 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(128 DOWNTO 128) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(64 DOWNTO 64)
									);
MUX_REORD_UPDATE_65 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(130 DOWNTO 130) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(65 DOWNTO 65)
									);
MUX_REORD_UPDATE_66 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(132 DOWNTO 132) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(66 DOWNTO 66)
									);
MUX_REORD_UPDATE_67 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(134 DOWNTO 134) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(67 DOWNTO 67)
									);
MUX_REORD_UPDATE_68 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(136 DOWNTO 136) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(68 DOWNTO 68)
									);
MUX_REORD_UPDATE_69 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(138 DOWNTO 138) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(69 DOWNTO 69)
									);
MUX_REORD_UPDATE_70 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(140 DOWNTO 140) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(70 DOWNTO 70)
									);
MUX_REORD_UPDATE_71 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(142 DOWNTO 142) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(71 DOWNTO 71)
									);
MUX_REORD_UPDATE_72 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(144 DOWNTO 144) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(72 DOWNTO 72)
									);
MUX_REORD_UPDATE_73 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(146 DOWNTO 146) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(73 DOWNTO 73)
									);
MUX_REORD_UPDATE_74 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(148 DOWNTO 148) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(74 DOWNTO 74)
									);
MUX_REORD_UPDATE_75 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(150 DOWNTO 150) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(75 DOWNTO 75)
									);
MUX_REORD_UPDATE_76 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(152 DOWNTO 152) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(76 DOWNTO 76)
									);
MUX_REORD_UPDATE_77 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(154 DOWNTO 154) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(77 DOWNTO 77)
									);
MUX_REORD_UPDATE_78 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(156 DOWNTO 156) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(78 DOWNTO 78)
									);
MUX_REORD_UPDATE_79 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(158 DOWNTO 158) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(79 DOWNTO 79)
									);
MUX_REORD_UPDATE_80 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(160 DOWNTO 160) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(80 DOWNTO 80)
									);
MUX_REORD_UPDATE_81 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(162 DOWNTO 162) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(81 DOWNTO 81)
									);
MUX_REORD_UPDATE_82 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(164 DOWNTO 164) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(82 DOWNTO 82)
									);
MUX_REORD_UPDATE_83 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(166 DOWNTO 166) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(83 DOWNTO 83)
									);
MUX_REORD_UPDATE_84 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(168 DOWNTO 168) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(84 DOWNTO 84)
									);
MUX_REORD_UPDATE_85 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(170 DOWNTO 170) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(85 DOWNTO 85)
									);
MUX_REORD_UPDATE_86 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(172 DOWNTO 172) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(86 DOWNTO 86)
									);
MUX_REORD_UPDATE_87 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(174 DOWNTO 174) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(87 DOWNTO 87)
									);
MUX_REORD_UPDATE_88 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(176 DOWNTO 176) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(88 DOWNTO 88)
									);
MUX_REORD_UPDATE_89 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(178 DOWNTO 178) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(89 DOWNTO 89)
									);
MUX_REORD_UPDATE_90 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(180 DOWNTO 180) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(90 DOWNTO 90)
									);
MUX_REORD_UPDATE_91 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(182 DOWNTO 182) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(91 DOWNTO 91)
									);
MUX_REORD_UPDATE_92 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(184 DOWNTO 184) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(92 DOWNTO 92)
									);
MUX_REORD_UPDATE_93 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(186 DOWNTO 186) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(93 DOWNTO 93)
									);
MUX_REORD_UPDATE_94 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(188 DOWNTO 188) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(94 DOWNTO 94)
									);
MUX_REORD_UPDATE_95 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(190 DOWNTO 190) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(95 DOWNTO 95)
									);
MUX_REORD_UPDATE_96 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(192 DOWNTO 192) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(96 DOWNTO 96)
									);
MUX_REORD_UPDATE_97 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(194 DOWNTO 194) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(97 DOWNTO 97)
									);
MUX_REORD_UPDATE_98 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(196 DOWNTO 196) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(98 DOWNTO 98)
									);
MUX_REORD_UPDATE_99 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(198 DOWNTO 198) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(99 DOWNTO 99)
									);
MUX_REORD_UPDATE_100 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(200 DOWNTO 200) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(100 DOWNTO 100)
									);
MUX_REORD_UPDATE_101 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(202 DOWNTO 202) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(101 DOWNTO 101)
									);
MUX_REORD_UPDATE_102 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(204 DOWNTO 204) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(102 DOWNTO 102)
									);
MUX_REORD_UPDATE_103 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(206 DOWNTO 206) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(103 DOWNTO 103)
									);
MUX_REORD_UPDATE_104 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(208 DOWNTO 208) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(104 DOWNTO 104)
									);
MUX_REORD_UPDATE_105 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(210 DOWNTO 210) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(105 DOWNTO 105)
									);
MUX_REORD_UPDATE_106 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(212 DOWNTO 212) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(106 DOWNTO 106)
									);
MUX_REORD_UPDATE_107 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(214 DOWNTO 214) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(107 DOWNTO 107)
									);
MUX_REORD_UPDATE_108 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(216 DOWNTO 216) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(108 DOWNTO 108)
									);
MUX_REORD_UPDATE_109 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(218 DOWNTO 218) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(109 DOWNTO 109)
									);
MUX_REORD_UPDATE_110 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(220 DOWNTO 220) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(110 DOWNTO 110)
									);
MUX_REORD_UPDATE_111 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(222 DOWNTO 222) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(111 DOWNTO 111)
									);
MUX_REORD_UPDATE_112 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(224 DOWNTO 224) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(112 DOWNTO 112)
									);
MUX_REORD_UPDATE_113 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(226 DOWNTO 226) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(113 DOWNTO 113)
									);
MUX_REORD_UPDATE_114 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(228 DOWNTO 228) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(114 DOWNTO 114)
									);
MUX_REORD_UPDATE_115 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(230 DOWNTO 230) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(115 DOWNTO 115)
									);
MUX_REORD_UPDATE_116 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(232 DOWNTO 232) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(116 DOWNTO 116)
									);
MUX_REORD_UPDATE_117 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(234 DOWNTO 234) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(117 DOWNTO 117)
									);
MUX_REORD_UPDATE_118 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(236 DOWNTO 236) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(118 DOWNTO 118)
									);
MUX_REORD_UPDATE_119 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(238 DOWNTO 238) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(119 DOWNTO 119)
									);
MUX_REORD_UPDATE_120 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(240 DOWNTO 240) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(120 DOWNTO 120)
									);
MUX_REORD_UPDATE_121 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(242 DOWNTO 242) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(121 DOWNTO 121)
									);
MUX_REORD_UPDATE_122 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(244 DOWNTO 244) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(122 DOWNTO 122)
									);
MUX_REORD_UPDATE_123 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(246 DOWNTO 246) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(123 DOWNTO 123)
									);
MUX_REORD_UPDATE_124 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(248 DOWNTO 248) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(124 DOWNTO 124)
									);
MUX_REORD_UPDATE_125 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(250 DOWNTO 250) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(125 DOWNTO 125)
									);
MUX_REORD_UPDATE_126 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(252 DOWNTO 252) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(126 DOWNTO 126)
									);
MUX_REORD_UPDATE_127 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(254 DOWNTO 254) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(127 DOWNTO 127)
									);
MUX_REORD_UPDATE_128 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(128 DOWNTO 128) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(256 DOWNTO 256) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(128 DOWNTO 128)
									);
MUX_REORD_UPDATE_129 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(258 DOWNTO 258) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(129 DOWNTO 129)
									);
MUX_REORD_UPDATE_130 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(130 DOWNTO 130) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(260 DOWNTO 260) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(130 DOWNTO 130)
									);
MUX_REORD_UPDATE_131 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(262 DOWNTO 262) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(131 DOWNTO 131)
									);
MUX_REORD_UPDATE_132 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(132 DOWNTO 132) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(264 DOWNTO 264) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(132 DOWNTO 132)
									);
MUX_REORD_UPDATE_133 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(266 DOWNTO 266) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(133 DOWNTO 133)
									);
MUX_REORD_UPDATE_134 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(134 DOWNTO 134) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(268 DOWNTO 268) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(134 DOWNTO 134)
									);
MUX_REORD_UPDATE_135 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(270 DOWNTO 270) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(135 DOWNTO 135)
									);
MUX_REORD_UPDATE_136 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(136 DOWNTO 136) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(272 DOWNTO 272) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(136 DOWNTO 136)
									);
MUX_REORD_UPDATE_137 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(274 DOWNTO 274) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(137 DOWNTO 137)
									);
MUX_REORD_UPDATE_138 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(138 DOWNTO 138) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(276 DOWNTO 276) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(138 DOWNTO 138)
									);
MUX_REORD_UPDATE_139 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(278 DOWNTO 278) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(139 DOWNTO 139)
									);
MUX_REORD_UPDATE_140 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(140 DOWNTO 140) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(280 DOWNTO 280) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(140 DOWNTO 140)
									);
MUX_REORD_UPDATE_141 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(282 DOWNTO 282) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(141 DOWNTO 141)
									);
MUX_REORD_UPDATE_142 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(142 DOWNTO 142) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(284 DOWNTO 284) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(142 DOWNTO 142)
									);
MUX_REORD_UPDATE_143 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(286 DOWNTO 286) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(143 DOWNTO 143)
									);
MUX_REORD_UPDATE_144 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(144 DOWNTO 144) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(288 DOWNTO 288) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(144 DOWNTO 144)
									);
MUX_REORD_UPDATE_145 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(290 DOWNTO 290) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(145 DOWNTO 145)
									);
MUX_REORD_UPDATE_146 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(146 DOWNTO 146) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(292 DOWNTO 292) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(146 DOWNTO 146)
									);
MUX_REORD_UPDATE_147 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(294 DOWNTO 294) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(147 DOWNTO 147)
									);
MUX_REORD_UPDATE_148 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(148 DOWNTO 148) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(296 DOWNTO 296) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(148 DOWNTO 148)
									);
MUX_REORD_UPDATE_149 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(298 DOWNTO 298) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(149 DOWNTO 149)
									);
MUX_REORD_UPDATE_150 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(150 DOWNTO 150) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(300 DOWNTO 300) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(150 DOWNTO 150)
									);
MUX_REORD_UPDATE_151 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(302 DOWNTO 302) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(151 DOWNTO 151)
									);
MUX_REORD_UPDATE_152 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(152 DOWNTO 152) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(304 DOWNTO 304) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(152 DOWNTO 152)
									);
MUX_REORD_UPDATE_153 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(306 DOWNTO 306) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(153 DOWNTO 153)
									);
MUX_REORD_UPDATE_154 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(154 DOWNTO 154) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(308 DOWNTO 308) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(154 DOWNTO 154)
									);
MUX_REORD_UPDATE_155 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(310 DOWNTO 310) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(155 DOWNTO 155)
									);
MUX_REORD_UPDATE_156 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(156 DOWNTO 156) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(312 DOWNTO 312) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(156 DOWNTO 156)
									);
MUX_REORD_UPDATE_157 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(314 DOWNTO 314) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(157 DOWNTO 157)
									);
MUX_REORD_UPDATE_158 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(158 DOWNTO 158) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(316 DOWNTO 316) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(158 DOWNTO 158)
									);
MUX_REORD_UPDATE_159 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(318 DOWNTO 318) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(159 DOWNTO 159)
									);
MUX_REORD_UPDATE_160 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(160 DOWNTO 160) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(320 DOWNTO 320) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(160 DOWNTO 160)
									);
MUX_REORD_UPDATE_161 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(322 DOWNTO 322) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(161 DOWNTO 161)
									);
MUX_REORD_UPDATE_162 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(162 DOWNTO 162) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(324 DOWNTO 324) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(162 DOWNTO 162)
									);
MUX_REORD_UPDATE_163 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(326 DOWNTO 326) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(163 DOWNTO 163)
									);
MUX_REORD_UPDATE_164 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(164 DOWNTO 164) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(328 DOWNTO 328) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(164 DOWNTO 164)
									);
MUX_REORD_UPDATE_165 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(330 DOWNTO 330) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(165 DOWNTO 165)
									);
MUX_REORD_UPDATE_166 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(166 DOWNTO 166) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(332 DOWNTO 332) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(166 DOWNTO 166)
									);
MUX_REORD_UPDATE_167 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(334 DOWNTO 334) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(167 DOWNTO 167)
									);
MUX_REORD_UPDATE_168 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(168 DOWNTO 168) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(336 DOWNTO 336) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(168 DOWNTO 168)
									);
MUX_REORD_UPDATE_169 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(338 DOWNTO 338) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(169 DOWNTO 169)
									);
MUX_REORD_UPDATE_170 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(170 DOWNTO 170) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(340 DOWNTO 340) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(170 DOWNTO 170)
									);
MUX_REORD_UPDATE_171 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(342 DOWNTO 342) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(171 DOWNTO 171)
									);
MUX_REORD_UPDATE_172 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(172 DOWNTO 172) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(344 DOWNTO 344) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(172 DOWNTO 172)
									);
MUX_REORD_UPDATE_173 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(346 DOWNTO 346) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(173 DOWNTO 173)
									);
MUX_REORD_UPDATE_174 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(174 DOWNTO 174) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(348 DOWNTO 348) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(174 DOWNTO 174)
									);
MUX_REORD_UPDATE_175 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(350 DOWNTO 350) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(175 DOWNTO 175)
									);
MUX_REORD_UPDATE_176 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(176 DOWNTO 176) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(352 DOWNTO 352) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(176 DOWNTO 176)
									);
MUX_REORD_UPDATE_177 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(354 DOWNTO 354) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(177 DOWNTO 177)
									);
MUX_REORD_UPDATE_178 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(178 DOWNTO 178) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(356 DOWNTO 356) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(178 DOWNTO 178)
									);
MUX_REORD_UPDATE_179 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(358 DOWNTO 358) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(179 DOWNTO 179)
									);
MUX_REORD_UPDATE_180 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(180 DOWNTO 180) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(360 DOWNTO 360) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(180 DOWNTO 180)
									);
MUX_REORD_UPDATE_181 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(362 DOWNTO 362) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(181 DOWNTO 181)
									);
MUX_REORD_UPDATE_182 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(182 DOWNTO 182) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(364 DOWNTO 364) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(182 DOWNTO 182)
									);
MUX_REORD_UPDATE_183 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(366 DOWNTO 366) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(183 DOWNTO 183)
									);
MUX_REORD_UPDATE_184 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(184 DOWNTO 184) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(368 DOWNTO 368) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(184 DOWNTO 184)
									);
MUX_REORD_UPDATE_185 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(370 DOWNTO 370) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(185 DOWNTO 185)
									);
MUX_REORD_UPDATE_186 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(186 DOWNTO 186) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(372 DOWNTO 372) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(186 DOWNTO 186)
									);
MUX_REORD_UPDATE_187 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(374 DOWNTO 374) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(187 DOWNTO 187)
									);
MUX_REORD_UPDATE_188 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(188 DOWNTO 188) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(376 DOWNTO 376) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(188 DOWNTO 188)
									);
MUX_REORD_UPDATE_189 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(378 DOWNTO 378) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(189 DOWNTO 189)
									);
MUX_REORD_UPDATE_190 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(190 DOWNTO 190) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(380 DOWNTO 380) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(190 DOWNTO 190)
									);
MUX_REORD_UPDATE_191 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(382 DOWNTO 382) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(191 DOWNTO 191)
									);
MUX_REORD_UPDATE_192 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(192 DOWNTO 192) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(384 DOWNTO 384) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(192 DOWNTO 192)
									);
MUX_REORD_UPDATE_193 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(386 DOWNTO 386) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(193 DOWNTO 193)
									);
MUX_REORD_UPDATE_194 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(194 DOWNTO 194) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(388 DOWNTO 388) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(194 DOWNTO 194)
									);
MUX_REORD_UPDATE_195 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(390 DOWNTO 390) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(195 DOWNTO 195)
									);
MUX_REORD_UPDATE_196 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(196 DOWNTO 196) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(392 DOWNTO 392) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(196 DOWNTO 196)
									);
MUX_REORD_UPDATE_197 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(394 DOWNTO 394) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(197 DOWNTO 197)
									);
MUX_REORD_UPDATE_198 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(198 DOWNTO 198) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(396 DOWNTO 396) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(198 DOWNTO 198)
									);
MUX_REORD_UPDATE_199 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(398 DOWNTO 398) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(199 DOWNTO 199)
									);
MUX_REORD_UPDATE_200 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(200 DOWNTO 200) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(400 DOWNTO 400) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(200 DOWNTO 200)
									);
MUX_REORD_UPDATE_201 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(402 DOWNTO 402) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(201 DOWNTO 201)
									);
MUX_REORD_UPDATE_202 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(202 DOWNTO 202) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(404 DOWNTO 404) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(202 DOWNTO 202)
									);
MUX_REORD_UPDATE_203 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(406 DOWNTO 406) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(203 DOWNTO 203)
									);
MUX_REORD_UPDATE_204 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(204 DOWNTO 204) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(408 DOWNTO 408) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(204 DOWNTO 204)
									);
MUX_REORD_UPDATE_205 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(410 DOWNTO 410) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(205 DOWNTO 205)
									);
MUX_REORD_UPDATE_206 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(206 DOWNTO 206) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(412 DOWNTO 412) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(206 DOWNTO 206)
									);
MUX_REORD_UPDATE_207 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(414 DOWNTO 414) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(207 DOWNTO 207)
									);
MUX_REORD_UPDATE_208 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(208 DOWNTO 208) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(416 DOWNTO 416) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(208 DOWNTO 208)
									);
MUX_REORD_UPDATE_209 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(418 DOWNTO 418) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(209 DOWNTO 209)
									);
MUX_REORD_UPDATE_210 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(210 DOWNTO 210) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(420 DOWNTO 420) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(210 DOWNTO 210)
									);
MUX_REORD_UPDATE_211 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(422 DOWNTO 422) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(211 DOWNTO 211)
									);
MUX_REORD_UPDATE_212 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(212 DOWNTO 212) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(424 DOWNTO 424) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(212 DOWNTO 212)
									);
MUX_REORD_UPDATE_213 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(426 DOWNTO 426) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(213 DOWNTO 213)
									);
MUX_REORD_UPDATE_214 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(214 DOWNTO 214) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(428 DOWNTO 428) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(214 DOWNTO 214)
									);
MUX_REORD_UPDATE_215 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(430 DOWNTO 430) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(215 DOWNTO 215)
									);
MUX_REORD_UPDATE_216 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(216 DOWNTO 216) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(432 DOWNTO 432) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(216 DOWNTO 216)
									);
MUX_REORD_UPDATE_217 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(434 DOWNTO 434) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(217 DOWNTO 217)
									);
MUX_REORD_UPDATE_218 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(218 DOWNTO 218) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(436 DOWNTO 436) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(218 DOWNTO 218)
									);
MUX_REORD_UPDATE_219 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(438 DOWNTO 438) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(219 DOWNTO 219)
									);
MUX_REORD_UPDATE_220 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(220 DOWNTO 220) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(440 DOWNTO 440) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(220 DOWNTO 220)
									);
MUX_REORD_UPDATE_221 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(442 DOWNTO 442) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(221 DOWNTO 221)
									);
MUX_REORD_UPDATE_222 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(222 DOWNTO 222) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(444 DOWNTO 444) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(222 DOWNTO 222)
									);
MUX_REORD_UPDATE_223 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(446 DOWNTO 446) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(223 DOWNTO 223)
									);
MUX_REORD_UPDATE_224 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(224 DOWNTO 224) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(448 DOWNTO 448) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(224 DOWNTO 224)
									);
MUX_REORD_UPDATE_225 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(450 DOWNTO 450) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(225 DOWNTO 225)
									);
MUX_REORD_UPDATE_226 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(226 DOWNTO 226) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(452 DOWNTO 452) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(226 DOWNTO 226)
									);
MUX_REORD_UPDATE_227 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(454 DOWNTO 454) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(227 DOWNTO 227)
									);
MUX_REORD_UPDATE_228 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(228 DOWNTO 228) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(456 DOWNTO 456) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(228 DOWNTO 228)
									);
MUX_REORD_UPDATE_229 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(458 DOWNTO 458) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(229 DOWNTO 229)
									);
MUX_REORD_UPDATE_230 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(230 DOWNTO 230) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(460 DOWNTO 460) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(230 DOWNTO 230)
									);
MUX_REORD_UPDATE_231 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(462 DOWNTO 462) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(231 DOWNTO 231)
									);
MUX_REORD_UPDATE_232 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(232 DOWNTO 232) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(464 DOWNTO 464) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(232 DOWNTO 232)
									);
MUX_REORD_UPDATE_233 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(466 DOWNTO 466) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(233 DOWNTO 233)
									);
MUX_REORD_UPDATE_234 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(234 DOWNTO 234) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(468 DOWNTO 468) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(234 DOWNTO 234)
									);
MUX_REORD_UPDATE_235 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(470 DOWNTO 470) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(235 DOWNTO 235)
									);
MUX_REORD_UPDATE_236 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(236 DOWNTO 236) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(472 DOWNTO 472) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(236 DOWNTO 236)
									);
MUX_REORD_UPDATE_237 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(474 DOWNTO 474) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(237 DOWNTO 237)
									);
MUX_REORD_UPDATE_238 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(238 DOWNTO 238) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(476 DOWNTO 476) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(238 DOWNTO 238)
									);
MUX_REORD_UPDATE_239 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(478 DOWNTO 478) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(239 DOWNTO 239)
									);
MUX_REORD_UPDATE_240 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(240 DOWNTO 240) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(480 DOWNTO 480) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(240 DOWNTO 240)
									);
MUX_REORD_UPDATE_241 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(482 DOWNTO 482) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(241 DOWNTO 241)
									);
MUX_REORD_UPDATE_242 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(242 DOWNTO 242) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(484 DOWNTO 484) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(242 DOWNTO 242)
									);
MUX_REORD_UPDATE_243 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(486 DOWNTO 486) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(243 DOWNTO 243)
									);
MUX_REORD_UPDATE_244 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(244 DOWNTO 244) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(488 DOWNTO 488) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(244 DOWNTO 244)
									);
MUX_REORD_UPDATE_245 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(490 DOWNTO 490) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(245 DOWNTO 245)
									);
MUX_REORD_UPDATE_246 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(246 DOWNTO 246) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(492 DOWNTO 492) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(246 DOWNTO 246)
									);
MUX_REORD_UPDATE_247 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(494 DOWNTO 494) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(247 DOWNTO 247)
									);
MUX_REORD_UPDATE_248 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(248 DOWNTO 248) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(496 DOWNTO 496) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(248 DOWNTO 248)
									);
MUX_REORD_UPDATE_249 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(498 DOWNTO 498) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(249 DOWNTO 249)
									);
MUX_REORD_UPDATE_250 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(250 DOWNTO 250) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(500 DOWNTO 500) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(250 DOWNTO 250)
									);
MUX_REORD_UPDATE_251 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(502 DOWNTO 502) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(251 DOWNTO 251)
									);
MUX_REORD_UPDATE_252 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(252 DOWNTO 252) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(504 DOWNTO 504) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(252 DOWNTO 252)
									);
MUX_REORD_UPDATE_253 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(506 DOWNTO 506) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(253 DOWNTO 253)
									);
MUX_REORD_UPDATE_254 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(254 DOWNTO 254) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(508 DOWNTO 508) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(254 DOWNTO 254)
									);
MUX_REORD_UPDATE_255 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(510 DOWNTO 510) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(255 DOWNTO 255)
									);
MUX_REORD_UPDATE_256 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(256 DOWNTO 256) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(512 DOWNTO 512) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(256 DOWNTO 256)
									);
MUX_REORD_UPDATE_257 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(514 DOWNTO 514) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(257 DOWNTO 257)
									);
MUX_REORD_UPDATE_258 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(258 DOWNTO 258) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(516 DOWNTO 516) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(258 DOWNTO 258)
									);
MUX_REORD_UPDATE_259 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(518 DOWNTO 518) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(259 DOWNTO 259)
									);
MUX_REORD_UPDATE_260 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(260 DOWNTO 260) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(520 DOWNTO 520) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(260 DOWNTO 260)
									);
MUX_REORD_UPDATE_261 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(522 DOWNTO 522) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(261 DOWNTO 261)
									);
MUX_REORD_UPDATE_262 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(262 DOWNTO 262) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(524 DOWNTO 524) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(262 DOWNTO 262)
									);
MUX_REORD_UPDATE_263 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(526 DOWNTO 526) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(263 DOWNTO 263)
									);
MUX_REORD_UPDATE_264 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(264 DOWNTO 264) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(528 DOWNTO 528) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(264 DOWNTO 264)
									);
MUX_REORD_UPDATE_265 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(530 DOWNTO 530) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(265 DOWNTO 265)
									);
MUX_REORD_UPDATE_266 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(266 DOWNTO 266) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(532 DOWNTO 532) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(266 DOWNTO 266)
									);
MUX_REORD_UPDATE_267 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(534 DOWNTO 534) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(267 DOWNTO 267)
									);
MUX_REORD_UPDATE_268 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(268 DOWNTO 268) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(536 DOWNTO 536) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(268 DOWNTO 268)
									);
MUX_REORD_UPDATE_269 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(538 DOWNTO 538) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(269 DOWNTO 269)
									);
MUX_REORD_UPDATE_270 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(270 DOWNTO 270) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(540 DOWNTO 540) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(270 DOWNTO 270)
									);
MUX_REORD_UPDATE_271 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(542 DOWNTO 542) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(271 DOWNTO 271)
									);
MUX_REORD_UPDATE_272 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(272 DOWNTO 272) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(544 DOWNTO 544) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(272 DOWNTO 272)
									);
MUX_REORD_UPDATE_273 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(546 DOWNTO 546) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(273 DOWNTO 273)
									);
MUX_REORD_UPDATE_274 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(274 DOWNTO 274) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(548 DOWNTO 548) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(274 DOWNTO 274)
									);
MUX_REORD_UPDATE_275 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(550 DOWNTO 550) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(275 DOWNTO 275)
									);
MUX_REORD_UPDATE_276 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(276 DOWNTO 276) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(552 DOWNTO 552) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(276 DOWNTO 276)
									);
MUX_REORD_UPDATE_277 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(554 DOWNTO 554) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(277 DOWNTO 277)
									);
MUX_REORD_UPDATE_278 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(278 DOWNTO 278) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(556 DOWNTO 556) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(278 DOWNTO 278)
									);
MUX_REORD_UPDATE_279 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(558 DOWNTO 558) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(279 DOWNTO 279)
									);
MUX_REORD_UPDATE_280 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(280 DOWNTO 280) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(560 DOWNTO 560) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(280 DOWNTO 280)
									);
MUX_REORD_UPDATE_281 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(562 DOWNTO 562) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(281 DOWNTO 281)
									);
MUX_REORD_UPDATE_282 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(282 DOWNTO 282) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(564 DOWNTO 564) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(282 DOWNTO 282)
									);
MUX_REORD_UPDATE_283 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(566 DOWNTO 566) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(283 DOWNTO 283)
									);
MUX_REORD_UPDATE_284 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(284 DOWNTO 284) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(568 DOWNTO 568) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(284 DOWNTO 284)
									);
MUX_REORD_UPDATE_285 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(570 DOWNTO 570) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(285 DOWNTO 285)
									);
MUX_REORD_UPDATE_286 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(286 DOWNTO 286) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(572 DOWNTO 572) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(286 DOWNTO 286)
									);
MUX_REORD_UPDATE_287 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(574 DOWNTO 574) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(287 DOWNTO 287)
									);
MUX_REORD_UPDATE_288 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(288 DOWNTO 288) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(576 DOWNTO 576) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(288 DOWNTO 288)
									);
MUX_REORD_UPDATE_289 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(578 DOWNTO 578) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(289 DOWNTO 289)
									);
MUX_REORD_UPDATE_290 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(290 DOWNTO 290) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(580 DOWNTO 580) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(290 DOWNTO 290)
									);
MUX_REORD_UPDATE_291 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(582 DOWNTO 582) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(291 DOWNTO 291)
									);
MUX_REORD_UPDATE_292 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(292 DOWNTO 292) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(584 DOWNTO 584) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(292 DOWNTO 292)
									);
MUX_REORD_UPDATE_293 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(586 DOWNTO 586) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(293 DOWNTO 293)
									);
MUX_REORD_UPDATE_294 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(294 DOWNTO 294) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(588 DOWNTO 588) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(294 DOWNTO 294)
									);
MUX_REORD_UPDATE_295 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(590 DOWNTO 590) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(295 DOWNTO 295)
									);
MUX_REORD_UPDATE_296 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(296 DOWNTO 296) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(592 DOWNTO 592) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(296 DOWNTO 296)
									);
MUX_REORD_UPDATE_297 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(594 DOWNTO 594) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(297 DOWNTO 297)
									);
MUX_REORD_UPDATE_298 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(298 DOWNTO 298) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(596 DOWNTO 596) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(298 DOWNTO 298)
									);
MUX_REORD_UPDATE_299 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(598 DOWNTO 598) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(299 DOWNTO 299)
									);
MUX_REORD_UPDATE_300 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(300 DOWNTO 300) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(600 DOWNTO 600) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(300 DOWNTO 300)
									);
MUX_REORD_UPDATE_301 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(602 DOWNTO 602) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(301 DOWNTO 301)
									);
MUX_REORD_UPDATE_302 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(302 DOWNTO 302) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(604 DOWNTO 604) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(302 DOWNTO 302)
									);
MUX_REORD_UPDATE_303 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(606 DOWNTO 606) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(303 DOWNTO 303)
									);
MUX_REORD_UPDATE_304 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(304 DOWNTO 304) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(608 DOWNTO 608) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(304 DOWNTO 304)
									);
MUX_REORD_UPDATE_305 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(610 DOWNTO 610) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(305 DOWNTO 305)
									);
MUX_REORD_UPDATE_306 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(306 DOWNTO 306) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(612 DOWNTO 612) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(306 DOWNTO 306)
									);
MUX_REORD_UPDATE_307 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(614 DOWNTO 614) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(307 DOWNTO 307)
									);
MUX_REORD_UPDATE_308 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(308 DOWNTO 308) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(616 DOWNTO 616) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(308 DOWNTO 308)
									);
MUX_REORD_UPDATE_309 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(618 DOWNTO 618) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(309 DOWNTO 309)
									);
MUX_REORD_UPDATE_310 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(310 DOWNTO 310) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(620 DOWNTO 620) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(310 DOWNTO 310)
									);
MUX_REORD_UPDATE_311 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(622 DOWNTO 622) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(311 DOWNTO 311)
									);
MUX_REORD_UPDATE_312 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(312 DOWNTO 312) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(624 DOWNTO 624) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(312 DOWNTO 312)
									);
MUX_REORD_UPDATE_313 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(626 DOWNTO 626) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(313 DOWNTO 313)
									);
MUX_REORD_UPDATE_314 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(314 DOWNTO 314) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(628 DOWNTO 628) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(314 DOWNTO 314)
									);
MUX_REORD_UPDATE_315 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(630 DOWNTO 630) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(315 DOWNTO 315)
									);
MUX_REORD_UPDATE_316 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(316 DOWNTO 316) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(632 DOWNTO 632) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(316 DOWNTO 316)
									);
MUX_REORD_UPDATE_317 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(634 DOWNTO 634) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(317 DOWNTO 317)
									);
MUX_REORD_UPDATE_318 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(318 DOWNTO 318) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(636 DOWNTO 636) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(318 DOWNTO 318)
									);
MUX_REORD_UPDATE_319 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(638 DOWNTO 638) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(319 DOWNTO 319)
									);
MUX_REORD_UPDATE_320 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(320 DOWNTO 320) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(129 DOWNTO 129) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(640 DOWNTO 640) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(320 DOWNTO 320)
									);
MUX_REORD_UPDATE_321 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(131 DOWNTO 131) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(642 DOWNTO 642) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(321 DOWNTO 321)
									);
MUX_REORD_UPDATE_322 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(322 DOWNTO 322) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(133 DOWNTO 133) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(644 DOWNTO 644) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(322 DOWNTO 322)
									);
MUX_REORD_UPDATE_323 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(135 DOWNTO 135) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(646 DOWNTO 646) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(323 DOWNTO 323)
									);
MUX_REORD_UPDATE_324 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(324 DOWNTO 324) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(137 DOWNTO 137) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(648 DOWNTO 648) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(324 DOWNTO 324)
									);
MUX_REORD_UPDATE_325 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(139 DOWNTO 139) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(650 DOWNTO 650) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(325 DOWNTO 325)
									);
MUX_REORD_UPDATE_326 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(326 DOWNTO 326) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(141 DOWNTO 141) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(652 DOWNTO 652) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(326 DOWNTO 326)
									);
MUX_REORD_UPDATE_327 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(143 DOWNTO 143) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(654 DOWNTO 654) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(327 DOWNTO 327)
									);
MUX_REORD_UPDATE_328 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(328 DOWNTO 328) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(145 DOWNTO 145) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(656 DOWNTO 656) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(328 DOWNTO 328)
									);
MUX_REORD_UPDATE_329 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(147 DOWNTO 147) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(658 DOWNTO 658) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(329 DOWNTO 329)
									);
MUX_REORD_UPDATE_330 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(330 DOWNTO 330) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(149 DOWNTO 149) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(660 DOWNTO 660) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(330 DOWNTO 330)
									);
MUX_REORD_UPDATE_331 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(151 DOWNTO 151) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(662 DOWNTO 662) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(331 DOWNTO 331)
									);
MUX_REORD_UPDATE_332 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(332 DOWNTO 332) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(153 DOWNTO 153) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(664 DOWNTO 664) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(332 DOWNTO 332)
									);
MUX_REORD_UPDATE_333 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(155 DOWNTO 155) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(666 DOWNTO 666) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(333 DOWNTO 333)
									);
MUX_REORD_UPDATE_334 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(334 DOWNTO 334) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(157 DOWNTO 157) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(668 DOWNTO 668) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(334 DOWNTO 334)
									);
MUX_REORD_UPDATE_335 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(159 DOWNTO 159) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(670 DOWNTO 670) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(335 DOWNTO 335)
									);
MUX_REORD_UPDATE_336 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(336 DOWNTO 336) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(161 DOWNTO 161) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(672 DOWNTO 672) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(336 DOWNTO 336)
									);
MUX_REORD_UPDATE_337 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(163 DOWNTO 163) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(674 DOWNTO 674) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(337 DOWNTO 337)
									);
MUX_REORD_UPDATE_338 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(338 DOWNTO 338) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(165 DOWNTO 165) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(676 DOWNTO 676) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(338 DOWNTO 338)
									);
MUX_REORD_UPDATE_339 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(167 DOWNTO 167) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(678 DOWNTO 678) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(339 DOWNTO 339)
									);
MUX_REORD_UPDATE_340 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(340 DOWNTO 340) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(169 DOWNTO 169) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(680 DOWNTO 680) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(340 DOWNTO 340)
									);
MUX_REORD_UPDATE_341 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(171 DOWNTO 171) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(682 DOWNTO 682) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(341 DOWNTO 341)
									);
MUX_REORD_UPDATE_342 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(342 DOWNTO 342) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(173 DOWNTO 173) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(684 DOWNTO 684) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(342 DOWNTO 342)
									);
MUX_REORD_UPDATE_343 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(175 DOWNTO 175) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(686 DOWNTO 686) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(343 DOWNTO 343)
									);
MUX_REORD_UPDATE_344 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(344 DOWNTO 344) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(177 DOWNTO 177) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(688 DOWNTO 688) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(344 DOWNTO 344)
									);
MUX_REORD_UPDATE_345 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(179 DOWNTO 179) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(690 DOWNTO 690) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(345 DOWNTO 345)
									);
MUX_REORD_UPDATE_346 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(346 DOWNTO 346) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(181 DOWNTO 181) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(692 DOWNTO 692) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(346 DOWNTO 346)
									);
MUX_REORD_UPDATE_347 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(183 DOWNTO 183) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(694 DOWNTO 694) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(347 DOWNTO 347)
									);
MUX_REORD_UPDATE_348 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(348 DOWNTO 348) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(185 DOWNTO 185) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(696 DOWNTO 696) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(348 DOWNTO 348)
									);
MUX_REORD_UPDATE_349 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(187 DOWNTO 187) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(698 DOWNTO 698) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(349 DOWNTO 349)
									);
MUX_REORD_UPDATE_350 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(350 DOWNTO 350) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(189 DOWNTO 189) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(700 DOWNTO 700) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(350 DOWNTO 350)
									);
MUX_REORD_UPDATE_351 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(191 DOWNTO 191) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(702 DOWNTO 702) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(351 DOWNTO 351)
									);
MUX_REORD_UPDATE_352 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(352 DOWNTO 352) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(193 DOWNTO 193) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(704 DOWNTO 704) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(352 DOWNTO 352)
									);
MUX_REORD_UPDATE_353 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(195 DOWNTO 195) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(706 DOWNTO 706) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(353 DOWNTO 353)
									);
MUX_REORD_UPDATE_354 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(354 DOWNTO 354) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(197 DOWNTO 197) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(708 DOWNTO 708) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(354 DOWNTO 354)
									);
MUX_REORD_UPDATE_355 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(199 DOWNTO 199) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(710 DOWNTO 710) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(355 DOWNTO 355)
									);
MUX_REORD_UPDATE_356 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(356 DOWNTO 356) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(201 DOWNTO 201) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(712 DOWNTO 712) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(356 DOWNTO 356)
									);
MUX_REORD_UPDATE_357 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(203 DOWNTO 203) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(714 DOWNTO 714) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(357 DOWNTO 357)
									);
MUX_REORD_UPDATE_358 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(358 DOWNTO 358) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(205 DOWNTO 205) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(716 DOWNTO 716) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(358 DOWNTO 358)
									);
MUX_REORD_UPDATE_359 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(207 DOWNTO 207) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(718 DOWNTO 718) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(359 DOWNTO 359)
									);
MUX_REORD_UPDATE_360 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(360 DOWNTO 360) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(209 DOWNTO 209) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(720 DOWNTO 720) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(360 DOWNTO 360)
									);
MUX_REORD_UPDATE_361 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(211 DOWNTO 211) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(722 DOWNTO 722) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(361 DOWNTO 361)
									);
MUX_REORD_UPDATE_362 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(362 DOWNTO 362) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(213 DOWNTO 213) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(724 DOWNTO 724) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(362 DOWNTO 362)
									);
MUX_REORD_UPDATE_363 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(215 DOWNTO 215) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(726 DOWNTO 726) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(363 DOWNTO 363)
									);
MUX_REORD_UPDATE_364 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(364 DOWNTO 364) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(217 DOWNTO 217) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(728 DOWNTO 728) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(364 DOWNTO 364)
									);
MUX_REORD_UPDATE_365 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(219 DOWNTO 219) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(730 DOWNTO 730) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(365 DOWNTO 365)
									);
MUX_REORD_UPDATE_366 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(366 DOWNTO 366) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(221 DOWNTO 221) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(732 DOWNTO 732) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(366 DOWNTO 366)
									);
MUX_REORD_UPDATE_367 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(223 DOWNTO 223) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(734 DOWNTO 734) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(367 DOWNTO 367)
									);
MUX_REORD_UPDATE_368 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(368 DOWNTO 368) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(225 DOWNTO 225) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(736 DOWNTO 736) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(368 DOWNTO 368)
									);
MUX_REORD_UPDATE_369 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(227 DOWNTO 227) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(738 DOWNTO 738) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(369 DOWNTO 369)
									);
MUX_REORD_UPDATE_370 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(370 DOWNTO 370) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(229 DOWNTO 229) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(740 DOWNTO 740) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(370 DOWNTO 370)
									);
MUX_REORD_UPDATE_371 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(231 DOWNTO 231) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(742 DOWNTO 742) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(371 DOWNTO 371)
									);
MUX_REORD_UPDATE_372 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(372 DOWNTO 372) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(233 DOWNTO 233) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(744 DOWNTO 744) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(372 DOWNTO 372)
									);
MUX_REORD_UPDATE_373 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(235 DOWNTO 235) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(746 DOWNTO 746) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(373 DOWNTO 373)
									);
MUX_REORD_UPDATE_374 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(374 DOWNTO 374) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(237 DOWNTO 237) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(748 DOWNTO 748) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(374 DOWNTO 374)
									);
MUX_REORD_UPDATE_375 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(239 DOWNTO 239) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(750 DOWNTO 750) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(375 DOWNTO 375)
									);
MUX_REORD_UPDATE_376 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(376 DOWNTO 376) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(241 DOWNTO 241) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(752 DOWNTO 752) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(376 DOWNTO 376)
									);
MUX_REORD_UPDATE_377 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(243 DOWNTO 243) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(754 DOWNTO 754) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(377 DOWNTO 377)
									);
MUX_REORD_UPDATE_378 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(378 DOWNTO 378) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(245 DOWNTO 245) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(756 DOWNTO 756) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(378 DOWNTO 378)
									);
MUX_REORD_UPDATE_379 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(247 DOWNTO 247) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(758 DOWNTO 758) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(379 DOWNTO 379)
									);
MUX_REORD_UPDATE_380 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(380 DOWNTO 380) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(249 DOWNTO 249) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(760 DOWNTO 760) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(380 DOWNTO 380)
									);
MUX_REORD_UPDATE_381 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(251 DOWNTO 251) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(762 DOWNTO 762) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(381 DOWNTO 381)
									);
MUX_REORD_UPDATE_382 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(382 DOWNTO 382) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(253 DOWNTO 253) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(764 DOWNTO 764) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(382 DOWNTO 382)
									);
MUX_REORD_UPDATE_383 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(255 DOWNTO 255) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(766 DOWNTO 766) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(383 DOWNTO 383)
									);
MUX_REORD_UPDATE_384 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(384 DOWNTO 384) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(257 DOWNTO 257) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(768 DOWNTO 768) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(384 DOWNTO 384)
									);
MUX_REORD_UPDATE_385 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(259 DOWNTO 259) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(770 DOWNTO 770) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(385 DOWNTO 385)
									);
MUX_REORD_UPDATE_386 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(386 DOWNTO 386) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(261 DOWNTO 261) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(772 DOWNTO 772) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(386 DOWNTO 386)
									);
MUX_REORD_UPDATE_387 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(263 DOWNTO 263) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(774 DOWNTO 774) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(387 DOWNTO 387)
									);
MUX_REORD_UPDATE_388 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(388 DOWNTO 388) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(265 DOWNTO 265) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(776 DOWNTO 776) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(388 DOWNTO 388)
									);
MUX_REORD_UPDATE_389 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(267 DOWNTO 267) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(778 DOWNTO 778) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(389 DOWNTO 389)
									);
MUX_REORD_UPDATE_390 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(390 DOWNTO 390) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(269 DOWNTO 269) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(780 DOWNTO 780) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(390 DOWNTO 390)
									);
MUX_REORD_UPDATE_391 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(271 DOWNTO 271) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(782 DOWNTO 782) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(391 DOWNTO 391)
									);
MUX_REORD_UPDATE_392 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(392 DOWNTO 392) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(273 DOWNTO 273) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(784 DOWNTO 784) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(392 DOWNTO 392)
									);
MUX_REORD_UPDATE_393 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(275 DOWNTO 275) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(786 DOWNTO 786) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(393 DOWNTO 393)
									);
MUX_REORD_UPDATE_394 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(394 DOWNTO 394) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(277 DOWNTO 277) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(788 DOWNTO 788) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(394 DOWNTO 394)
									);
MUX_REORD_UPDATE_395 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(279 DOWNTO 279) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(790 DOWNTO 790) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(395 DOWNTO 395)
									);
MUX_REORD_UPDATE_396 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(396 DOWNTO 396) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(281 DOWNTO 281) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(792 DOWNTO 792) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(396 DOWNTO 396)
									);
MUX_REORD_UPDATE_397 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(283 DOWNTO 283) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(794 DOWNTO 794) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(397 DOWNTO 397)
									);
MUX_REORD_UPDATE_398 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(398 DOWNTO 398) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(285 DOWNTO 285) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(796 DOWNTO 796) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(398 DOWNTO 398)
									);
MUX_REORD_UPDATE_399 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(287 DOWNTO 287) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(798 DOWNTO 798) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(399 DOWNTO 399)
									);
MUX_REORD_UPDATE_400 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(400 DOWNTO 400) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(289 DOWNTO 289) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(800 DOWNTO 800) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(400 DOWNTO 400)
									);
MUX_REORD_UPDATE_401 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(291 DOWNTO 291) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(802 DOWNTO 802) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(401 DOWNTO 401)
									);
MUX_REORD_UPDATE_402 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(402 DOWNTO 402) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(293 DOWNTO 293) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(804 DOWNTO 804) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(402 DOWNTO 402)
									);
MUX_REORD_UPDATE_403 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(295 DOWNTO 295) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(806 DOWNTO 806) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(403 DOWNTO 403)
									);
MUX_REORD_UPDATE_404 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(404 DOWNTO 404) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(297 DOWNTO 297) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(808 DOWNTO 808) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(404 DOWNTO 404)
									);
MUX_REORD_UPDATE_405 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(299 DOWNTO 299) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(810 DOWNTO 810) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(405 DOWNTO 405)
									);
MUX_REORD_UPDATE_406 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(406 DOWNTO 406) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(301 DOWNTO 301) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(812 DOWNTO 812) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(406 DOWNTO 406)
									);
MUX_REORD_UPDATE_407 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(303 DOWNTO 303) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(814 DOWNTO 814) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(407 DOWNTO 407)
									);
MUX_REORD_UPDATE_408 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(408 DOWNTO 408) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(305 DOWNTO 305) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(816 DOWNTO 816) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(408 DOWNTO 408)
									);
MUX_REORD_UPDATE_409 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(307 DOWNTO 307) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(818 DOWNTO 818) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(409 DOWNTO 409)
									);
MUX_REORD_UPDATE_410 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(410 DOWNTO 410) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(309 DOWNTO 309) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(820 DOWNTO 820) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(410 DOWNTO 410)
									);
MUX_REORD_UPDATE_411 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(311 DOWNTO 311) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(822 DOWNTO 822) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(411 DOWNTO 411)
									);
MUX_REORD_UPDATE_412 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(412 DOWNTO 412) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(313 DOWNTO 313) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(824 DOWNTO 824) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(412 DOWNTO 412)
									);
MUX_REORD_UPDATE_413 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(315 DOWNTO 315) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(826 DOWNTO 826) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(413 DOWNTO 413)
									);
MUX_REORD_UPDATE_414 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(414 DOWNTO 414) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(317 DOWNTO 317) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(828 DOWNTO 828) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(414 DOWNTO 414)
									);
MUX_REORD_UPDATE_415 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(319 DOWNTO 319) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(830 DOWNTO 830) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(415 DOWNTO 415)
									);
MUX_REORD_UPDATE_416 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(416 DOWNTO 416) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(321 DOWNTO 321) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(832 DOWNTO 832) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(416 DOWNTO 416)
									);
MUX_REORD_UPDATE_417 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(323 DOWNTO 323) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(834 DOWNTO 834) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(417 DOWNTO 417)
									);
MUX_REORD_UPDATE_418 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(418 DOWNTO 418) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(325 DOWNTO 325) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(836 DOWNTO 836) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(418 DOWNTO 418)
									);
MUX_REORD_UPDATE_419 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(327 DOWNTO 327) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(838 DOWNTO 838) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(419 DOWNTO 419)
									);
MUX_REORD_UPDATE_420 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(420 DOWNTO 420) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(329 DOWNTO 329) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(840 DOWNTO 840) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(420 DOWNTO 420)
									);
MUX_REORD_UPDATE_421 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(331 DOWNTO 331) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(842 DOWNTO 842) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(421 DOWNTO 421)
									);
MUX_REORD_UPDATE_422 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(422 DOWNTO 422) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(333 DOWNTO 333) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(844 DOWNTO 844) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(422 DOWNTO 422)
									);
MUX_REORD_UPDATE_423 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(335 DOWNTO 335) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(846 DOWNTO 846) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(423 DOWNTO 423)
									);
MUX_REORD_UPDATE_424 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(424 DOWNTO 424) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(337 DOWNTO 337) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(848 DOWNTO 848) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(424 DOWNTO 424)
									);
MUX_REORD_UPDATE_425 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(339 DOWNTO 339) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(850 DOWNTO 850) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(425 DOWNTO 425)
									);
MUX_REORD_UPDATE_426 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(426 DOWNTO 426) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(341 DOWNTO 341) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(852 DOWNTO 852) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(426 DOWNTO 426)
									);
MUX_REORD_UPDATE_427 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(343 DOWNTO 343) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(854 DOWNTO 854) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(427 DOWNTO 427)
									);
MUX_REORD_UPDATE_428 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(428 DOWNTO 428) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(345 DOWNTO 345) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(856 DOWNTO 856) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(428 DOWNTO 428)
									);
MUX_REORD_UPDATE_429 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(347 DOWNTO 347) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(858 DOWNTO 858) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(429 DOWNTO 429)
									);
MUX_REORD_UPDATE_430 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(430 DOWNTO 430) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(349 DOWNTO 349) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(860 DOWNTO 860) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(430 DOWNTO 430)
									);
MUX_REORD_UPDATE_431 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(351 DOWNTO 351) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(862 DOWNTO 862) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(431 DOWNTO 431)
									);
MUX_REORD_UPDATE_432 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(432 DOWNTO 432) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(353 DOWNTO 353) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(864 DOWNTO 864) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(432 DOWNTO 432)
									);
MUX_REORD_UPDATE_433 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(355 DOWNTO 355) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(866 DOWNTO 866) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(433 DOWNTO 433)
									);
MUX_REORD_UPDATE_434 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(434 DOWNTO 434) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(357 DOWNTO 357) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(868 DOWNTO 868) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(434 DOWNTO 434)
									);
MUX_REORD_UPDATE_435 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(359 DOWNTO 359) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(870 DOWNTO 870) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(435 DOWNTO 435)
									);
MUX_REORD_UPDATE_436 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(436 DOWNTO 436) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(361 DOWNTO 361) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(872 DOWNTO 872) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(436 DOWNTO 436)
									);
MUX_REORD_UPDATE_437 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(363 DOWNTO 363) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(874 DOWNTO 874) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(437 DOWNTO 437)
									);
MUX_REORD_UPDATE_438 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(438 DOWNTO 438) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(365 DOWNTO 365) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(876 DOWNTO 876) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(438 DOWNTO 438)
									);
MUX_REORD_UPDATE_439 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(367 DOWNTO 367) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(878 DOWNTO 878) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(439 DOWNTO 439)
									);
MUX_REORD_UPDATE_440 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(440 DOWNTO 440) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(369 DOWNTO 369) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(880 DOWNTO 880) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(440 DOWNTO 440)
									);
MUX_REORD_UPDATE_441 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(371 DOWNTO 371) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(882 DOWNTO 882) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(441 DOWNTO 441)
									);
MUX_REORD_UPDATE_442 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(442 DOWNTO 442) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(373 DOWNTO 373) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(884 DOWNTO 884) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(442 DOWNTO 442)
									);
MUX_REORD_UPDATE_443 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(375 DOWNTO 375) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(886 DOWNTO 886) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(443 DOWNTO 443)
									);
MUX_REORD_UPDATE_444 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(444 DOWNTO 444) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(377 DOWNTO 377) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(888 DOWNTO 888) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(444 DOWNTO 444)
									);
MUX_REORD_UPDATE_445 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(379 DOWNTO 379) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(890 DOWNTO 890) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(445 DOWNTO 445)
									);
MUX_REORD_UPDATE_446 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(446 DOWNTO 446) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(381 DOWNTO 381) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(892 DOWNTO 892) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(446 DOWNTO 446)
									);
MUX_REORD_UPDATE_447 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(383 DOWNTO 383) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(894 DOWNTO 894) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(447 DOWNTO 447)
									);
MUX_REORD_UPDATE_448 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(448 DOWNTO 448) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(385 DOWNTO 385) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(896 DOWNTO 896) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(448 DOWNTO 448)
									);
MUX_REORD_UPDATE_449 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(387 DOWNTO 387) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(898 DOWNTO 898) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(449 DOWNTO 449)
									);
MUX_REORD_UPDATE_450 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(450 DOWNTO 450) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(389 DOWNTO 389) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(900 DOWNTO 900) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(450 DOWNTO 450)
									);
MUX_REORD_UPDATE_451 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(391 DOWNTO 391) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(902 DOWNTO 902) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(451 DOWNTO 451)
									);
MUX_REORD_UPDATE_452 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(452 DOWNTO 452) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(393 DOWNTO 393) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(904 DOWNTO 904) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(452 DOWNTO 452)
									);
MUX_REORD_UPDATE_453 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(395 DOWNTO 395) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(906 DOWNTO 906) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(453 DOWNTO 453)
									);
MUX_REORD_UPDATE_454 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(454 DOWNTO 454) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(397 DOWNTO 397) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(908 DOWNTO 908) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(454 DOWNTO 454)
									);
MUX_REORD_UPDATE_455 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(399 DOWNTO 399) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(910 DOWNTO 910) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(455 DOWNTO 455)
									);
MUX_REORD_UPDATE_456 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(456 DOWNTO 456) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(401 DOWNTO 401) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(912 DOWNTO 912) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(456 DOWNTO 456)
									);
MUX_REORD_UPDATE_457 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(403 DOWNTO 403) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(914 DOWNTO 914) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(457 DOWNTO 457)
									);
MUX_REORD_UPDATE_458 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(458 DOWNTO 458) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(405 DOWNTO 405) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(916 DOWNTO 916) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(458 DOWNTO 458)
									);
MUX_REORD_UPDATE_459 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(407 DOWNTO 407) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(918 DOWNTO 918) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(459 DOWNTO 459)
									);
MUX_REORD_UPDATE_460 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(460 DOWNTO 460) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(409 DOWNTO 409) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(920 DOWNTO 920) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(460 DOWNTO 460)
									);
MUX_REORD_UPDATE_461 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(411 DOWNTO 411) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(922 DOWNTO 922) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(461 DOWNTO 461)
									);
MUX_REORD_UPDATE_462 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(462 DOWNTO 462) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(413 DOWNTO 413) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(924 DOWNTO 924) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(462 DOWNTO 462)
									);
MUX_REORD_UPDATE_463 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(415 DOWNTO 415) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(926 DOWNTO 926) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(463 DOWNTO 463)
									);
MUX_REORD_UPDATE_464 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(464 DOWNTO 464) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(417 DOWNTO 417) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(928 DOWNTO 928) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(464 DOWNTO 464)
									);
MUX_REORD_UPDATE_465 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(419 DOWNTO 419) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(930 DOWNTO 930) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(465 DOWNTO 465)
									);
MUX_REORD_UPDATE_466 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(466 DOWNTO 466) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(421 DOWNTO 421) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(932 DOWNTO 932) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(466 DOWNTO 466)
									);
MUX_REORD_UPDATE_467 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(423 DOWNTO 423) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(934 DOWNTO 934) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(467 DOWNTO 467)
									);
MUX_REORD_UPDATE_468 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(468 DOWNTO 468) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(425 DOWNTO 425) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(936 DOWNTO 936) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(468 DOWNTO 468)
									);
MUX_REORD_UPDATE_469 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(427 DOWNTO 427) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(938 DOWNTO 938) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(469 DOWNTO 469)
									);
MUX_REORD_UPDATE_470 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(470 DOWNTO 470) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(429 DOWNTO 429) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(940 DOWNTO 940) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(470 DOWNTO 470)
									);
MUX_REORD_UPDATE_471 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(431 DOWNTO 431) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(942 DOWNTO 942) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(471 DOWNTO 471)
									);
MUX_REORD_UPDATE_472 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(472 DOWNTO 472) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(433 DOWNTO 433) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(944 DOWNTO 944) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(472 DOWNTO 472)
									);
MUX_REORD_UPDATE_473 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(435 DOWNTO 435) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(946 DOWNTO 946) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(473 DOWNTO 473)
									);
MUX_REORD_UPDATE_474 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(474 DOWNTO 474) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(437 DOWNTO 437) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(948 DOWNTO 948) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(474 DOWNTO 474)
									);
MUX_REORD_UPDATE_475 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(439 DOWNTO 439) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(950 DOWNTO 950) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(475 DOWNTO 475)
									);
MUX_REORD_UPDATE_476 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(476 DOWNTO 476) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(441 DOWNTO 441) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(952 DOWNTO 952) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(476 DOWNTO 476)
									);
MUX_REORD_UPDATE_477 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(443 DOWNTO 443) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(954 DOWNTO 954) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(477 DOWNTO 477)
									);
MUX_REORD_UPDATE_478 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(478 DOWNTO 478) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(445 DOWNTO 445) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(956 DOWNTO 956) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(478 DOWNTO 478)
									);
MUX_REORD_UPDATE_479 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(447 DOWNTO 447) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(958 DOWNTO 958) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(479 DOWNTO 479)
									);
MUX_REORD_UPDATE_480 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(480 DOWNTO 480) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(449 DOWNTO 449) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(960 DOWNTO 960) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(480 DOWNTO 480)
									);
MUX_REORD_UPDATE_481 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(451 DOWNTO 451) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(962 DOWNTO 962) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(481 DOWNTO 481)
									);
MUX_REORD_UPDATE_482 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(482 DOWNTO 482) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(453 DOWNTO 453) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(964 DOWNTO 964) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(482 DOWNTO 482)
									);
MUX_REORD_UPDATE_483 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(455 DOWNTO 455) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(966 DOWNTO 966) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(483 DOWNTO 483)
									);
MUX_REORD_UPDATE_484 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(484 DOWNTO 484) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(457 DOWNTO 457) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(968 DOWNTO 968) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(484 DOWNTO 484)
									);
MUX_REORD_UPDATE_485 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(459 DOWNTO 459) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(970 DOWNTO 970) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(485 DOWNTO 485)
									);
MUX_REORD_UPDATE_486 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(486 DOWNTO 486) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(461 DOWNTO 461) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(972 DOWNTO 972) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(486 DOWNTO 486)
									);
MUX_REORD_UPDATE_487 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(463 DOWNTO 463) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(974 DOWNTO 974) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(487 DOWNTO 487)
									);
MUX_REORD_UPDATE_488 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(488 DOWNTO 488) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(465 DOWNTO 465) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(976 DOWNTO 976) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(488 DOWNTO 488)
									);
MUX_REORD_UPDATE_489 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(467 DOWNTO 467) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(978 DOWNTO 978) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(489 DOWNTO 489)
									);
MUX_REORD_UPDATE_490 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(490 DOWNTO 490) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(469 DOWNTO 469) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(980 DOWNTO 980) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(490 DOWNTO 490)
									);
MUX_REORD_UPDATE_491 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(471 DOWNTO 471) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(982 DOWNTO 982) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(491 DOWNTO 491)
									);
MUX_REORD_UPDATE_492 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(492 DOWNTO 492) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(473 DOWNTO 473) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(984 DOWNTO 984) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(492 DOWNTO 492)
									);
MUX_REORD_UPDATE_493 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(475 DOWNTO 475) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(986 DOWNTO 986) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(493 DOWNTO 493)
									);
MUX_REORD_UPDATE_494 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(494 DOWNTO 494) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(477 DOWNTO 477) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(988 DOWNTO 988) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(494 DOWNTO 494)
									);
MUX_REORD_UPDATE_495 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(479 DOWNTO 479) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(990 DOWNTO 990) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(495 DOWNTO 495)
									);
MUX_REORD_UPDATE_496 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(496 DOWNTO 496) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(481 DOWNTO 481) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(992 DOWNTO 992) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(496 DOWNTO 496)
									);
MUX_REORD_UPDATE_497 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(483 DOWNTO 483) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(994 DOWNTO 994) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(497 DOWNTO 497)
									);
MUX_REORD_UPDATE_498 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(498 DOWNTO 498) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(485 DOWNTO 485) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(996 DOWNTO 996) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(498 DOWNTO 498)
									);
MUX_REORD_UPDATE_499 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(487 DOWNTO 487) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(998 DOWNTO 998) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(499 DOWNTO 499)
									);
MUX_REORD_UPDATE_500 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(500 DOWNTO 500) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(489 DOWNTO 489) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(500 DOWNTO 500)
									);
MUX_REORD_UPDATE_501 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(491 DOWNTO 491) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(501 DOWNTO 501)
									);
MUX_REORD_UPDATE_502 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(502 DOWNTO 502) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(493 DOWNTO 493) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(502 DOWNTO 502)
									);
MUX_REORD_UPDATE_503 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(495 DOWNTO 495) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(503 DOWNTO 503)
									);
MUX_REORD_UPDATE_504 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(504 DOWNTO 504) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(497 DOWNTO 497) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(504 DOWNTO 504)
									);
MUX_REORD_UPDATE_505 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(499 DOWNTO 499) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(505 DOWNTO 505)
									);
MUX_REORD_UPDATE_506 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(506 DOWNTO 506) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(501 DOWNTO 501) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(506 DOWNTO 506)
									);
MUX_REORD_UPDATE_507 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(503 DOWNTO 503) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(507 DOWNTO 507)
									);
MUX_REORD_UPDATE_508 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(508 DOWNTO 508) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(505 DOWNTO 505) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(508 DOWNTO 508)
									);
MUX_REORD_UPDATE_509 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(507 DOWNTO 507) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(509 DOWNTO 509)
									);
MUX_REORD_UPDATE_510 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(510 DOWNTO 510) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(509 DOWNTO 509) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(510 DOWNTO 510)
									);
MUX_REORD_UPDATE_511 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(511 DOWNTO 511) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(511 DOWNTO 511)
									);
MUX_REORD_UPDATE_512 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(512 DOWNTO 512) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1 DOWNTO 1) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(512 DOWNTO 512)
									);
MUX_REORD_UPDATE_513 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(3 DOWNTO 3) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(513 DOWNTO 513)
									);
MUX_REORD_UPDATE_514 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(514 DOWNTO 514) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(5 DOWNTO 5) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(514 DOWNTO 514)
									);
MUX_REORD_UPDATE_515 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(7 DOWNTO 7) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(515 DOWNTO 515)
									);
MUX_REORD_UPDATE_516 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(516 DOWNTO 516) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(9 DOWNTO 9) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(516 DOWNTO 516)
									);
MUX_REORD_UPDATE_517 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(11 DOWNTO 11) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(517 DOWNTO 517)
									);
MUX_REORD_UPDATE_518 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(518 DOWNTO 518) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(13 DOWNTO 13) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(518 DOWNTO 518)
									);
MUX_REORD_UPDATE_519 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(15 DOWNTO 15) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(519 DOWNTO 519)
									);
MUX_REORD_UPDATE_520 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(520 DOWNTO 520) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(17 DOWNTO 17) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(520 DOWNTO 520)
									);
MUX_REORD_UPDATE_521 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(19 DOWNTO 19) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(521 DOWNTO 521)
									);
MUX_REORD_UPDATE_522 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(522 DOWNTO 522) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(21 DOWNTO 21) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(522 DOWNTO 522)
									);
MUX_REORD_UPDATE_523 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(23 DOWNTO 23) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(523 DOWNTO 523)
									);
MUX_REORD_UPDATE_524 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(524 DOWNTO 524) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(25 DOWNTO 25) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(524 DOWNTO 524)
									);
MUX_REORD_UPDATE_525 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(27 DOWNTO 27) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(525 DOWNTO 525)
									);
MUX_REORD_UPDATE_526 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(526 DOWNTO 526) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(29 DOWNTO 29) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(526 DOWNTO 526)
									);
MUX_REORD_UPDATE_527 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(31 DOWNTO 31) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(527 DOWNTO 527)
									);
MUX_REORD_UPDATE_528 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(528 DOWNTO 528) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(33 DOWNTO 33) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(528 DOWNTO 528)
									);
MUX_REORD_UPDATE_529 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(35 DOWNTO 35) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(529 DOWNTO 529)
									);
MUX_REORD_UPDATE_530 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(530 DOWNTO 530) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(37 DOWNTO 37) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(530 DOWNTO 530)
									);
MUX_REORD_UPDATE_531 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(39 DOWNTO 39) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(531 DOWNTO 531)
									);
MUX_REORD_UPDATE_532 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(532 DOWNTO 532) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(41 DOWNTO 41) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(532 DOWNTO 532)
									);
MUX_REORD_UPDATE_533 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(43 DOWNTO 43) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(533 DOWNTO 533)
									);
MUX_REORD_UPDATE_534 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(534 DOWNTO 534) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(45 DOWNTO 45) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(534 DOWNTO 534)
									);
MUX_REORD_UPDATE_535 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(47 DOWNTO 47) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(535 DOWNTO 535)
									);
MUX_REORD_UPDATE_536 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(536 DOWNTO 536) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(49 DOWNTO 49) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(536 DOWNTO 536)
									);
MUX_REORD_UPDATE_537 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(51 DOWNTO 51) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(537 DOWNTO 537)
									);
MUX_REORD_UPDATE_538 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(538 DOWNTO 538) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(53 DOWNTO 53) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(538 DOWNTO 538)
									);
MUX_REORD_UPDATE_539 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(55 DOWNTO 55) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(539 DOWNTO 539)
									);
MUX_REORD_UPDATE_540 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(540 DOWNTO 540) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(57 DOWNTO 57) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(540 DOWNTO 540)
									);
MUX_REORD_UPDATE_541 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(59 DOWNTO 59) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(541 DOWNTO 541)
									);
MUX_REORD_UPDATE_542 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(542 DOWNTO 542) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(61 DOWNTO 61) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(542 DOWNTO 542)
									);
MUX_REORD_UPDATE_543 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(63 DOWNTO 63) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(543 DOWNTO 543)
									);
MUX_REORD_UPDATE_544 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(544 DOWNTO 544) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(65 DOWNTO 65) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(544 DOWNTO 544)
									);
MUX_REORD_UPDATE_545 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(67 DOWNTO 67) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(545 DOWNTO 545)
									);
MUX_REORD_UPDATE_546 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(546 DOWNTO 546) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(69 DOWNTO 69) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(546 DOWNTO 546)
									);
MUX_REORD_UPDATE_547 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(71 DOWNTO 71) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(547 DOWNTO 547)
									);
MUX_REORD_UPDATE_548 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(548 DOWNTO 548) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(73 DOWNTO 73) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(548 DOWNTO 548)
									);
MUX_REORD_UPDATE_549 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(75 DOWNTO 75) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(549 DOWNTO 549)
									);
MUX_REORD_UPDATE_550 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(550 DOWNTO 550) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(77 DOWNTO 77) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(550 DOWNTO 550)
									);
MUX_REORD_UPDATE_551 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(79 DOWNTO 79) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(551 DOWNTO 551)
									);
MUX_REORD_UPDATE_552 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(552 DOWNTO 552) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(81 DOWNTO 81) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(552 DOWNTO 552)
									);
MUX_REORD_UPDATE_553 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(83 DOWNTO 83) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(553 DOWNTO 553)
									);
MUX_REORD_UPDATE_554 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(554 DOWNTO 554) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(85 DOWNTO 85) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(554 DOWNTO 554)
									);
MUX_REORD_UPDATE_555 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(87 DOWNTO 87) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(555 DOWNTO 555)
									);
MUX_REORD_UPDATE_556 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(556 DOWNTO 556) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(89 DOWNTO 89) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(556 DOWNTO 556)
									);
MUX_REORD_UPDATE_557 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(91 DOWNTO 91) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(557 DOWNTO 557)
									);
MUX_REORD_UPDATE_558 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(558 DOWNTO 558) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(93 DOWNTO 93) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(558 DOWNTO 558)
									);
MUX_REORD_UPDATE_559 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(95 DOWNTO 95) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(559 DOWNTO 559)
									);
MUX_REORD_UPDATE_560 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(560 DOWNTO 560) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(97 DOWNTO 97) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(560 DOWNTO 560)
									);
MUX_REORD_UPDATE_561 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(99 DOWNTO 99) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(561 DOWNTO 561)
									);
MUX_REORD_UPDATE_562 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(562 DOWNTO 562) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(101 DOWNTO 101) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(562 DOWNTO 562)
									);
MUX_REORD_UPDATE_563 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(103 DOWNTO 103) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(563 DOWNTO 563)
									);
MUX_REORD_UPDATE_564 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(564 DOWNTO 564) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(105 DOWNTO 105) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(564 DOWNTO 564)
									);
MUX_REORD_UPDATE_565 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(107 DOWNTO 107) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(565 DOWNTO 565)
									);
MUX_REORD_UPDATE_566 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(566 DOWNTO 566) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(109 DOWNTO 109) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(566 DOWNTO 566)
									);
MUX_REORD_UPDATE_567 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(111 DOWNTO 111) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(567 DOWNTO 567)
									);
MUX_REORD_UPDATE_568 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(568 DOWNTO 568) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(113 DOWNTO 113) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(568 DOWNTO 568)
									);
MUX_REORD_UPDATE_569 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(115 DOWNTO 115) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(569 DOWNTO 569)
									);
MUX_REORD_UPDATE_570 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(570 DOWNTO 570) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(117 DOWNTO 117) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(570 DOWNTO 570)
									);
MUX_REORD_UPDATE_571 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(119 DOWNTO 119) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(571 DOWNTO 571)
									);
MUX_REORD_UPDATE_572 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(572 DOWNTO 572) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(121 DOWNTO 121) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(572 DOWNTO 572)
									);
MUX_REORD_UPDATE_573 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(123 DOWNTO 123) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(573 DOWNTO 573)
									);
MUX_REORD_UPDATE_574 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(574 DOWNTO 574) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(125 DOWNTO 125) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(574 DOWNTO 574)
									);
MUX_REORD_UPDATE_575 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(127 DOWNTO 127) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(575 DOWNTO 575)
									);
MUX_REORD_UPDATE_576 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(576 DOWNTO 576) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(129 DOWNTO 129) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(576 DOWNTO 576)
									);
MUX_REORD_UPDATE_577 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(131 DOWNTO 131) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(577 DOWNTO 577)
									);
MUX_REORD_UPDATE_578 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(578 DOWNTO 578) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(133 DOWNTO 133) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(578 DOWNTO 578)
									);
MUX_REORD_UPDATE_579 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(135 DOWNTO 135) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(579 DOWNTO 579)
									);
MUX_REORD_UPDATE_580 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(580 DOWNTO 580) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(137 DOWNTO 137) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(580 DOWNTO 580)
									);
MUX_REORD_UPDATE_581 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(139 DOWNTO 139) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(581 DOWNTO 581)
									);
MUX_REORD_UPDATE_582 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(582 DOWNTO 582) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(141 DOWNTO 141) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(582 DOWNTO 582)
									);
MUX_REORD_UPDATE_583 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(143 DOWNTO 143) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(583 DOWNTO 583)
									);
MUX_REORD_UPDATE_584 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(584 DOWNTO 584) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(145 DOWNTO 145) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(584 DOWNTO 584)
									);
MUX_REORD_UPDATE_585 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(147 DOWNTO 147) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(585 DOWNTO 585)
									);
MUX_REORD_UPDATE_586 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(586 DOWNTO 586) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(149 DOWNTO 149) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(586 DOWNTO 586)
									);
MUX_REORD_UPDATE_587 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(151 DOWNTO 151) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(587 DOWNTO 587)
									);
MUX_REORD_UPDATE_588 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(588 DOWNTO 588) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(153 DOWNTO 153) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(588 DOWNTO 588)
									);
MUX_REORD_UPDATE_589 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(155 DOWNTO 155) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(589 DOWNTO 589)
									);
MUX_REORD_UPDATE_590 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(590 DOWNTO 590) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(157 DOWNTO 157) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(590 DOWNTO 590)
									);
MUX_REORD_UPDATE_591 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(159 DOWNTO 159) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(591 DOWNTO 591)
									);
MUX_REORD_UPDATE_592 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(592 DOWNTO 592) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(161 DOWNTO 161) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(592 DOWNTO 592)
									);
MUX_REORD_UPDATE_593 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(163 DOWNTO 163) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(593 DOWNTO 593)
									);
MUX_REORD_UPDATE_594 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(594 DOWNTO 594) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(165 DOWNTO 165) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(594 DOWNTO 594)
									);
MUX_REORD_UPDATE_595 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(167 DOWNTO 167) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(595 DOWNTO 595)
									);
MUX_REORD_UPDATE_596 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(596 DOWNTO 596) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(169 DOWNTO 169) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(596 DOWNTO 596)
									);
MUX_REORD_UPDATE_597 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(171 DOWNTO 171) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(597 DOWNTO 597)
									);
MUX_REORD_UPDATE_598 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(598 DOWNTO 598) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(173 DOWNTO 173) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(598 DOWNTO 598)
									);
MUX_REORD_UPDATE_599 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(175 DOWNTO 175) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(599 DOWNTO 599)
									);
MUX_REORD_UPDATE_600 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(600 DOWNTO 600) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(177 DOWNTO 177) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(600 DOWNTO 600)
									);
MUX_REORD_UPDATE_601 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(179 DOWNTO 179) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(601 DOWNTO 601)
									);
MUX_REORD_UPDATE_602 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(602 DOWNTO 602) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(181 DOWNTO 181) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(602 DOWNTO 602)
									);
MUX_REORD_UPDATE_603 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(183 DOWNTO 183) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(603 DOWNTO 603)
									);
MUX_REORD_UPDATE_604 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(604 DOWNTO 604) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(185 DOWNTO 185) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(604 DOWNTO 604)
									);
MUX_REORD_UPDATE_605 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(187 DOWNTO 187) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(605 DOWNTO 605)
									);
MUX_REORD_UPDATE_606 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(606 DOWNTO 606) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(189 DOWNTO 189) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(606 DOWNTO 606)
									);
MUX_REORD_UPDATE_607 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(191 DOWNTO 191) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(607 DOWNTO 607)
									);
MUX_REORD_UPDATE_608 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(608 DOWNTO 608) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(193 DOWNTO 193) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(608 DOWNTO 608)
									);
MUX_REORD_UPDATE_609 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(195 DOWNTO 195) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(609 DOWNTO 609)
									);
MUX_REORD_UPDATE_610 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(610 DOWNTO 610) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(197 DOWNTO 197) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(610 DOWNTO 610)
									);
MUX_REORD_UPDATE_611 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(199 DOWNTO 199) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(611 DOWNTO 611)
									);
MUX_REORD_UPDATE_612 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(612 DOWNTO 612) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(201 DOWNTO 201) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(612 DOWNTO 612)
									);
MUX_REORD_UPDATE_613 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(203 DOWNTO 203) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(613 DOWNTO 613)
									);
MUX_REORD_UPDATE_614 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(614 DOWNTO 614) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(205 DOWNTO 205) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(614 DOWNTO 614)
									);
MUX_REORD_UPDATE_615 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(207 DOWNTO 207) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(615 DOWNTO 615)
									);
MUX_REORD_UPDATE_616 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(616 DOWNTO 616) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(209 DOWNTO 209) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(616 DOWNTO 616)
									);
MUX_REORD_UPDATE_617 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(211 DOWNTO 211) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(617 DOWNTO 617)
									);
MUX_REORD_UPDATE_618 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(618 DOWNTO 618) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(213 DOWNTO 213) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(618 DOWNTO 618)
									);
MUX_REORD_UPDATE_619 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(215 DOWNTO 215) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(619 DOWNTO 619)
									);
MUX_REORD_UPDATE_620 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(620 DOWNTO 620) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(217 DOWNTO 217) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(620 DOWNTO 620)
									);
MUX_REORD_UPDATE_621 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(219 DOWNTO 219) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(621 DOWNTO 621)
									);
MUX_REORD_UPDATE_622 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(622 DOWNTO 622) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(221 DOWNTO 221) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(622 DOWNTO 622)
									);
MUX_REORD_UPDATE_623 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(223 DOWNTO 223) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(623 DOWNTO 623)
									);
MUX_REORD_UPDATE_624 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(624 DOWNTO 624) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(225 DOWNTO 225) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(624 DOWNTO 624)
									);
MUX_REORD_UPDATE_625 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(227 DOWNTO 227) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(625 DOWNTO 625)
									);
MUX_REORD_UPDATE_626 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(626 DOWNTO 626) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(229 DOWNTO 229) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(626 DOWNTO 626)
									);
MUX_REORD_UPDATE_627 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(231 DOWNTO 231) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(627 DOWNTO 627)
									);
MUX_REORD_UPDATE_628 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(628 DOWNTO 628) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(233 DOWNTO 233) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(628 DOWNTO 628)
									);
MUX_REORD_UPDATE_629 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(235 DOWNTO 235) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(629 DOWNTO 629)
									);
MUX_REORD_UPDATE_630 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(630 DOWNTO 630) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(237 DOWNTO 237) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(630 DOWNTO 630)
									);
MUX_REORD_UPDATE_631 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(239 DOWNTO 239) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(631 DOWNTO 631)
									);
MUX_REORD_UPDATE_632 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(632 DOWNTO 632) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(241 DOWNTO 241) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(632 DOWNTO 632)
									);
MUX_REORD_UPDATE_633 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(243 DOWNTO 243) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(633 DOWNTO 633)
									);
MUX_REORD_UPDATE_634 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(634 DOWNTO 634) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(245 DOWNTO 245) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(634 DOWNTO 634)
									);
MUX_REORD_UPDATE_635 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(247 DOWNTO 247) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(635 DOWNTO 635)
									);
MUX_REORD_UPDATE_636 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(636 DOWNTO 636) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(249 DOWNTO 249) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(636 DOWNTO 636)
									);
MUX_REORD_UPDATE_637 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(251 DOWNTO 251) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(637 DOWNTO 637)
									);
MUX_REORD_UPDATE_638 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(638 DOWNTO 638) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(253 DOWNTO 253) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(638 DOWNTO 638)
									);
MUX_REORD_UPDATE_639 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(255 DOWNTO 255) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(639 DOWNTO 639)
									);
MUX_REORD_UPDATE_640 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(640 DOWNTO 640) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(257 DOWNTO 257) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(640 DOWNTO 640)
									);
MUX_REORD_UPDATE_641 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(259 DOWNTO 259) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(641 DOWNTO 641)
									);
MUX_REORD_UPDATE_642 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(642 DOWNTO 642) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(261 DOWNTO 261) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(642 DOWNTO 642)
									);
MUX_REORD_UPDATE_643 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(263 DOWNTO 263) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(643 DOWNTO 643)
									);
MUX_REORD_UPDATE_644 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(644 DOWNTO 644) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(265 DOWNTO 265) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(644 DOWNTO 644)
									);
MUX_REORD_UPDATE_645 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(267 DOWNTO 267) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(645 DOWNTO 645)
									);
MUX_REORD_UPDATE_646 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(646 DOWNTO 646) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(269 DOWNTO 269) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(646 DOWNTO 646)
									);
MUX_REORD_UPDATE_647 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(271 DOWNTO 271) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(647 DOWNTO 647)
									);
MUX_REORD_UPDATE_648 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(648 DOWNTO 648) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(273 DOWNTO 273) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(648 DOWNTO 648)
									);
MUX_REORD_UPDATE_649 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(275 DOWNTO 275) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(649 DOWNTO 649)
									);
MUX_REORD_UPDATE_650 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(650 DOWNTO 650) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(277 DOWNTO 277) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(650 DOWNTO 650)
									);
MUX_REORD_UPDATE_651 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(279 DOWNTO 279) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(651 DOWNTO 651)
									);
MUX_REORD_UPDATE_652 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(652 DOWNTO 652) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(281 DOWNTO 281) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(652 DOWNTO 652)
									);
MUX_REORD_UPDATE_653 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(283 DOWNTO 283) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(653 DOWNTO 653)
									);
MUX_REORD_UPDATE_654 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(654 DOWNTO 654) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(285 DOWNTO 285) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(654 DOWNTO 654)
									);
MUX_REORD_UPDATE_655 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(287 DOWNTO 287) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(655 DOWNTO 655)
									);
MUX_REORD_UPDATE_656 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(656 DOWNTO 656) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(289 DOWNTO 289) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(656 DOWNTO 656)
									);
MUX_REORD_UPDATE_657 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(291 DOWNTO 291) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(657 DOWNTO 657)
									);
MUX_REORD_UPDATE_658 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(658 DOWNTO 658) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(293 DOWNTO 293) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(658 DOWNTO 658)
									);
MUX_REORD_UPDATE_659 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(295 DOWNTO 295) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(659 DOWNTO 659)
									);
MUX_REORD_UPDATE_660 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(660 DOWNTO 660) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(297 DOWNTO 297) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(660 DOWNTO 660)
									);
MUX_REORD_UPDATE_661 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(299 DOWNTO 299) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(661 DOWNTO 661)
									);
MUX_REORD_UPDATE_662 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(662 DOWNTO 662) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(301 DOWNTO 301) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(662 DOWNTO 662)
									);
MUX_REORD_UPDATE_663 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(303 DOWNTO 303) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(663 DOWNTO 663)
									);
MUX_REORD_UPDATE_664 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(664 DOWNTO 664) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(305 DOWNTO 305) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(664 DOWNTO 664)
									);
MUX_REORD_UPDATE_665 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(307 DOWNTO 307) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(665 DOWNTO 665)
									);
MUX_REORD_UPDATE_666 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(666 DOWNTO 666) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(309 DOWNTO 309) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(666 DOWNTO 666)
									);
MUX_REORD_UPDATE_667 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(311 DOWNTO 311) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(667 DOWNTO 667)
									);
MUX_REORD_UPDATE_668 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(668 DOWNTO 668) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(313 DOWNTO 313) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(668 DOWNTO 668)
									);
MUX_REORD_UPDATE_669 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(315 DOWNTO 315) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(669 DOWNTO 669)
									);
MUX_REORD_UPDATE_670 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(670 DOWNTO 670) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(317 DOWNTO 317) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(670 DOWNTO 670)
									);
MUX_REORD_UPDATE_671 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(319 DOWNTO 319) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(671 DOWNTO 671)
									);
MUX_REORD_UPDATE_672 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(672 DOWNTO 672) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(321 DOWNTO 321) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(672 DOWNTO 672)
									);
MUX_REORD_UPDATE_673 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(323 DOWNTO 323) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(673 DOWNTO 673)
									);
MUX_REORD_UPDATE_674 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(674 DOWNTO 674) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(325 DOWNTO 325) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(674 DOWNTO 674)
									);
MUX_REORD_UPDATE_675 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(327 DOWNTO 327) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(675 DOWNTO 675)
									);
MUX_REORD_UPDATE_676 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(676 DOWNTO 676) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(329 DOWNTO 329) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(676 DOWNTO 676)
									);
MUX_REORD_UPDATE_677 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(331 DOWNTO 331) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(677 DOWNTO 677)
									);
MUX_REORD_UPDATE_678 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(678 DOWNTO 678) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(333 DOWNTO 333) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(678 DOWNTO 678)
									);
MUX_REORD_UPDATE_679 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(335 DOWNTO 335) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(679 DOWNTO 679)
									);
MUX_REORD_UPDATE_680 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(680 DOWNTO 680) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(337 DOWNTO 337) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(680 DOWNTO 680)
									);
MUX_REORD_UPDATE_681 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(339 DOWNTO 339) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(681 DOWNTO 681)
									);
MUX_REORD_UPDATE_682 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(682 DOWNTO 682) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(341 DOWNTO 341) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(682 DOWNTO 682)
									);
MUX_REORD_UPDATE_683 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(343 DOWNTO 343) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(683 DOWNTO 683)
									);
MUX_REORD_UPDATE_684 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(684 DOWNTO 684) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(345 DOWNTO 345) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(684 DOWNTO 684)
									);
MUX_REORD_UPDATE_685 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(347 DOWNTO 347) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(685 DOWNTO 685)
									);
MUX_REORD_UPDATE_686 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(686 DOWNTO 686) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(349 DOWNTO 349) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(686 DOWNTO 686)
									);
MUX_REORD_UPDATE_687 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(351 DOWNTO 351) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(687 DOWNTO 687)
									);
MUX_REORD_UPDATE_688 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(688 DOWNTO 688) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(353 DOWNTO 353) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(688 DOWNTO 688)
									);
MUX_REORD_UPDATE_689 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(355 DOWNTO 355) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(689 DOWNTO 689)
									);
MUX_REORD_UPDATE_690 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(690 DOWNTO 690) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(357 DOWNTO 357) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(690 DOWNTO 690)
									);
MUX_REORD_UPDATE_691 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(359 DOWNTO 359) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(691 DOWNTO 691)
									);
MUX_REORD_UPDATE_692 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(692 DOWNTO 692) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(361 DOWNTO 361) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(692 DOWNTO 692)
									);
MUX_REORD_UPDATE_693 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(363 DOWNTO 363) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(693 DOWNTO 693)
									);
MUX_REORD_UPDATE_694 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(694 DOWNTO 694) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(365 DOWNTO 365) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(694 DOWNTO 694)
									);
MUX_REORD_UPDATE_695 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(367 DOWNTO 367) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(695 DOWNTO 695)
									);
MUX_REORD_UPDATE_696 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(696 DOWNTO 696) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(369 DOWNTO 369) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(696 DOWNTO 696)
									);
MUX_REORD_UPDATE_697 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(371 DOWNTO 371) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(697 DOWNTO 697)
									);
MUX_REORD_UPDATE_698 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(698 DOWNTO 698) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(373 DOWNTO 373) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(698 DOWNTO 698)
									);
MUX_REORD_UPDATE_699 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(375 DOWNTO 375) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(699 DOWNTO 699)
									);
MUX_REORD_UPDATE_700 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(700 DOWNTO 700) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(377 DOWNTO 377) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(700 DOWNTO 700)
									);
MUX_REORD_UPDATE_701 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(379 DOWNTO 379) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(701 DOWNTO 701)
									);
MUX_REORD_UPDATE_702 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(702 DOWNTO 702) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(381 DOWNTO 381) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(702 DOWNTO 702)
									);
MUX_REORD_UPDATE_703 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(383 DOWNTO 383) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(703 DOWNTO 703)
									);
MUX_REORD_UPDATE_704 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(704 DOWNTO 704) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(385 DOWNTO 385) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(704 DOWNTO 704)
									);
MUX_REORD_UPDATE_705 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(387 DOWNTO 387) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(705 DOWNTO 705)
									);
MUX_REORD_UPDATE_706 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(706 DOWNTO 706) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(389 DOWNTO 389) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(706 DOWNTO 706)
									);
MUX_REORD_UPDATE_707 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(391 DOWNTO 391) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(707 DOWNTO 707)
									);
MUX_REORD_UPDATE_708 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(708 DOWNTO 708) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(393 DOWNTO 393) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(708 DOWNTO 708)
									);
MUX_REORD_UPDATE_709 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(395 DOWNTO 395) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(709 DOWNTO 709)
									);
MUX_REORD_UPDATE_710 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(710 DOWNTO 710) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(397 DOWNTO 397) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(710 DOWNTO 710)
									);
MUX_REORD_UPDATE_711 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(399 DOWNTO 399) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(711 DOWNTO 711)
									);
MUX_REORD_UPDATE_712 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(712 DOWNTO 712) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(401 DOWNTO 401) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(712 DOWNTO 712)
									);
MUX_REORD_UPDATE_713 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(403 DOWNTO 403) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(713 DOWNTO 713)
									);
MUX_REORD_UPDATE_714 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(714 DOWNTO 714) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(405 DOWNTO 405) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(714 DOWNTO 714)
									);
MUX_REORD_UPDATE_715 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(407 DOWNTO 407) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(715 DOWNTO 715)
									);
MUX_REORD_UPDATE_716 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(716 DOWNTO 716) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(409 DOWNTO 409) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(716 DOWNTO 716)
									);
MUX_REORD_UPDATE_717 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(411 DOWNTO 411) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(717 DOWNTO 717)
									);
MUX_REORD_UPDATE_718 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(718 DOWNTO 718) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(413 DOWNTO 413) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(718 DOWNTO 718)
									);
MUX_REORD_UPDATE_719 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(415 DOWNTO 415) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(719 DOWNTO 719)
									);
MUX_REORD_UPDATE_720 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(720 DOWNTO 720) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(417 DOWNTO 417) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(720 DOWNTO 720)
									);
MUX_REORD_UPDATE_721 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(419 DOWNTO 419) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(721 DOWNTO 721)
									);
MUX_REORD_UPDATE_722 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(722 DOWNTO 722) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(421 DOWNTO 421) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(722 DOWNTO 722)
									);
MUX_REORD_UPDATE_723 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(423 DOWNTO 423) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(723 DOWNTO 723)
									);
MUX_REORD_UPDATE_724 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(724 DOWNTO 724) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(425 DOWNTO 425) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(724 DOWNTO 724)
									);
MUX_REORD_UPDATE_725 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(427 DOWNTO 427) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(725 DOWNTO 725)
									);
MUX_REORD_UPDATE_726 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(726 DOWNTO 726) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(429 DOWNTO 429) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(726 DOWNTO 726)
									);
MUX_REORD_UPDATE_727 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(431 DOWNTO 431) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(727 DOWNTO 727)
									);
MUX_REORD_UPDATE_728 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(728 DOWNTO 728) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(433 DOWNTO 433) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(728 DOWNTO 728)
									);
MUX_REORD_UPDATE_729 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(435 DOWNTO 435) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(729 DOWNTO 729)
									);
MUX_REORD_UPDATE_730 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(730 DOWNTO 730) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(437 DOWNTO 437) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(730 DOWNTO 730)
									);
MUX_REORD_UPDATE_731 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(439 DOWNTO 439) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(731 DOWNTO 731)
									);
MUX_REORD_UPDATE_732 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(732 DOWNTO 732) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(441 DOWNTO 441) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(732 DOWNTO 732)
									);
MUX_REORD_UPDATE_733 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(443 DOWNTO 443) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(733 DOWNTO 733)
									);
MUX_REORD_UPDATE_734 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(734 DOWNTO 734) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(445 DOWNTO 445) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(734 DOWNTO 734)
									);
MUX_REORD_UPDATE_735 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(447 DOWNTO 447) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(735 DOWNTO 735)
									);
MUX_REORD_UPDATE_736 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(736 DOWNTO 736) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(449 DOWNTO 449) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(736 DOWNTO 736)
									);
MUX_REORD_UPDATE_737 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(451 DOWNTO 451) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(737 DOWNTO 737)
									);
MUX_REORD_UPDATE_738 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(738 DOWNTO 738) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(453 DOWNTO 453) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(738 DOWNTO 738)
									);
MUX_REORD_UPDATE_739 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(455 DOWNTO 455) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(739 DOWNTO 739)
									);
MUX_REORD_UPDATE_740 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(740 DOWNTO 740) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(457 DOWNTO 457) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(740 DOWNTO 740)
									);
MUX_REORD_UPDATE_741 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(459 DOWNTO 459) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(741 DOWNTO 741)
									);
MUX_REORD_UPDATE_742 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(742 DOWNTO 742) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(461 DOWNTO 461) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(742 DOWNTO 742)
									);
MUX_REORD_UPDATE_743 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(463 DOWNTO 463) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(743 DOWNTO 743)
									);
MUX_REORD_UPDATE_744 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(744 DOWNTO 744) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(465 DOWNTO 465) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(744 DOWNTO 744)
									);
MUX_REORD_UPDATE_745 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(467 DOWNTO 467) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(745 DOWNTO 745)
									);
MUX_REORD_UPDATE_746 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(746 DOWNTO 746) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(469 DOWNTO 469) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(746 DOWNTO 746)
									);
MUX_REORD_UPDATE_747 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(471 DOWNTO 471) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(747 DOWNTO 747)
									);
MUX_REORD_UPDATE_748 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(748 DOWNTO 748) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(473 DOWNTO 473) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(748 DOWNTO 748)
									);
MUX_REORD_UPDATE_749 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(475 DOWNTO 475) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(749 DOWNTO 749)
									);
MUX_REORD_UPDATE_750 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(750 DOWNTO 750) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(477 DOWNTO 477) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(750 DOWNTO 750)
									);
MUX_REORD_UPDATE_751 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(479 DOWNTO 479) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(751 DOWNTO 751)
									);
MUX_REORD_UPDATE_752 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(752 DOWNTO 752) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(481 DOWNTO 481) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(752 DOWNTO 752)
									);
MUX_REORD_UPDATE_753 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(483 DOWNTO 483) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(753 DOWNTO 753)
									);
MUX_REORD_UPDATE_754 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(754 DOWNTO 754) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(485 DOWNTO 485) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(754 DOWNTO 754)
									);
MUX_REORD_UPDATE_755 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(487 DOWNTO 487) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(755 DOWNTO 755)
									);
MUX_REORD_UPDATE_756 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(756 DOWNTO 756) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(489 DOWNTO 489) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(756 DOWNTO 756)
									);
MUX_REORD_UPDATE_757 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(491 DOWNTO 491) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(757 DOWNTO 757)
									);
MUX_REORD_UPDATE_758 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(758 DOWNTO 758) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(493 DOWNTO 493) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(758 DOWNTO 758)
									);
MUX_REORD_UPDATE_759 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(495 DOWNTO 495) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(759 DOWNTO 759)
									);
MUX_REORD_UPDATE_760 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(760 DOWNTO 760) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(497 DOWNTO 497) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(760 DOWNTO 760)
									);
MUX_REORD_UPDATE_761 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(499 DOWNTO 499) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(761 DOWNTO 761)
									);
MUX_REORD_UPDATE_762 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(762 DOWNTO 762) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(501 DOWNTO 501) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(762 DOWNTO 762)
									);
MUX_REORD_UPDATE_763 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(503 DOWNTO 503) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(763 DOWNTO 763)
									);
MUX_REORD_UPDATE_764 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(764 DOWNTO 764) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(505 DOWNTO 505) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(764 DOWNTO 764)
									);
MUX_REORD_UPDATE_765 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(507 DOWNTO 507) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(765 DOWNTO 765)
									);
MUX_REORD_UPDATE_766 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(766 DOWNTO 766) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(509 DOWNTO 509) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(766 DOWNTO 766)
									);
MUX_REORD_UPDATE_767 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(511 DOWNTO 511) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(767 DOWNTO 767)
									);
MUX_REORD_UPDATE_768 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(768 DOWNTO 768) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(513 DOWNTO 513) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(513 DOWNTO 513) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(768 DOWNTO 768)
									);
MUX_REORD_UPDATE_769 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(515 DOWNTO 515) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(515 DOWNTO 515) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(769 DOWNTO 769)
									);
MUX_REORD_UPDATE_770 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(770 DOWNTO 770) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(517 DOWNTO 517) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(517 DOWNTO 517) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(770 DOWNTO 770)
									);
MUX_REORD_UPDATE_771 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(519 DOWNTO 519) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(519 DOWNTO 519) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(771 DOWNTO 771)
									);
MUX_REORD_UPDATE_772 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(772 DOWNTO 772) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(521 DOWNTO 521) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(521 DOWNTO 521) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(772 DOWNTO 772)
									);
MUX_REORD_UPDATE_773 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(523 DOWNTO 523) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(523 DOWNTO 523) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(773 DOWNTO 773)
									);
MUX_REORD_UPDATE_774 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(774 DOWNTO 774) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(525 DOWNTO 525) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(525 DOWNTO 525) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(774 DOWNTO 774)
									);
MUX_REORD_UPDATE_775 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(527 DOWNTO 527) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(527 DOWNTO 527) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(775 DOWNTO 775)
									);
MUX_REORD_UPDATE_776 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(776 DOWNTO 776) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(529 DOWNTO 529) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(529 DOWNTO 529) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(776 DOWNTO 776)
									);
MUX_REORD_UPDATE_777 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(531 DOWNTO 531) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(531 DOWNTO 531) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(777 DOWNTO 777)
									);
MUX_REORD_UPDATE_778 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(778 DOWNTO 778) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(533 DOWNTO 533) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(533 DOWNTO 533) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(778 DOWNTO 778)
									);
MUX_REORD_UPDATE_779 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(535 DOWNTO 535) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(535 DOWNTO 535) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(779 DOWNTO 779)
									);
MUX_REORD_UPDATE_780 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(780 DOWNTO 780) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(537 DOWNTO 537) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(537 DOWNTO 537) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(780 DOWNTO 780)
									);
MUX_REORD_UPDATE_781 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(539 DOWNTO 539) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(539 DOWNTO 539) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(781 DOWNTO 781)
									);
MUX_REORD_UPDATE_782 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(782 DOWNTO 782) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(541 DOWNTO 541) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(541 DOWNTO 541) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(782 DOWNTO 782)
									);
MUX_REORD_UPDATE_783 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(543 DOWNTO 543) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(543 DOWNTO 543) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(783 DOWNTO 783)
									);
MUX_REORD_UPDATE_784 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(784 DOWNTO 784) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(545 DOWNTO 545) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(545 DOWNTO 545) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(784 DOWNTO 784)
									);
MUX_REORD_UPDATE_785 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(547 DOWNTO 547) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(547 DOWNTO 547) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(785 DOWNTO 785)
									);
MUX_REORD_UPDATE_786 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(786 DOWNTO 786) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(549 DOWNTO 549) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(549 DOWNTO 549) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(786 DOWNTO 786)
									);
MUX_REORD_UPDATE_787 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(551 DOWNTO 551) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(551 DOWNTO 551) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(787 DOWNTO 787)
									);
MUX_REORD_UPDATE_788 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(788 DOWNTO 788) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(553 DOWNTO 553) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(553 DOWNTO 553) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(788 DOWNTO 788)
									);
MUX_REORD_UPDATE_789 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(555 DOWNTO 555) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(555 DOWNTO 555) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(789 DOWNTO 789)
									);
MUX_REORD_UPDATE_790 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(790 DOWNTO 790) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(557 DOWNTO 557) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(557 DOWNTO 557) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(790 DOWNTO 790)
									);
MUX_REORD_UPDATE_791 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(559 DOWNTO 559) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(559 DOWNTO 559) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(791 DOWNTO 791)
									);
MUX_REORD_UPDATE_792 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(792 DOWNTO 792) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(561 DOWNTO 561) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(561 DOWNTO 561) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(792 DOWNTO 792)
									);
MUX_REORD_UPDATE_793 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(563 DOWNTO 563) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(563 DOWNTO 563) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(793 DOWNTO 793)
									);
MUX_REORD_UPDATE_794 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(794 DOWNTO 794) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(565 DOWNTO 565) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(565 DOWNTO 565) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(794 DOWNTO 794)
									);
MUX_REORD_UPDATE_795 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(567 DOWNTO 567) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(567 DOWNTO 567) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(795 DOWNTO 795)
									);
MUX_REORD_UPDATE_796 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(796 DOWNTO 796) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(569 DOWNTO 569) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(569 DOWNTO 569) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(796 DOWNTO 796)
									);
MUX_REORD_UPDATE_797 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(571 DOWNTO 571) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(571 DOWNTO 571) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(797 DOWNTO 797)
									);
MUX_REORD_UPDATE_798 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(798 DOWNTO 798) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(573 DOWNTO 573) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(573 DOWNTO 573) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(798 DOWNTO 798)
									);
MUX_REORD_UPDATE_799 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(575 DOWNTO 575) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(575 DOWNTO 575) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(799 DOWNTO 799)
									);
MUX_REORD_UPDATE_800 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(800 DOWNTO 800) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(577 DOWNTO 577) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(577 DOWNTO 577) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(800 DOWNTO 800)
									);
MUX_REORD_UPDATE_801 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(579 DOWNTO 579) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(579 DOWNTO 579) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(801 DOWNTO 801)
									);
MUX_REORD_UPDATE_802 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(802 DOWNTO 802) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(581 DOWNTO 581) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(581 DOWNTO 581) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(802 DOWNTO 802)
									);
MUX_REORD_UPDATE_803 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(583 DOWNTO 583) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(583 DOWNTO 583) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(803 DOWNTO 803)
									);
MUX_REORD_UPDATE_804 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(804 DOWNTO 804) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(585 DOWNTO 585) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(585 DOWNTO 585) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(804 DOWNTO 804)
									);
MUX_REORD_UPDATE_805 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(587 DOWNTO 587) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(587 DOWNTO 587) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(805 DOWNTO 805)
									);
MUX_REORD_UPDATE_806 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(806 DOWNTO 806) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(589 DOWNTO 589) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(589 DOWNTO 589) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(806 DOWNTO 806)
									);
MUX_REORD_UPDATE_807 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(591 DOWNTO 591) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(591 DOWNTO 591) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(807 DOWNTO 807)
									);
MUX_REORD_UPDATE_808 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(808 DOWNTO 808) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(593 DOWNTO 593) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(593 DOWNTO 593) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(808 DOWNTO 808)
									);
MUX_REORD_UPDATE_809 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(595 DOWNTO 595) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(595 DOWNTO 595) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(809 DOWNTO 809)
									);
MUX_REORD_UPDATE_810 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(810 DOWNTO 810) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(597 DOWNTO 597) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(597 DOWNTO 597) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(810 DOWNTO 810)
									);
MUX_REORD_UPDATE_811 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(599 DOWNTO 599) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(599 DOWNTO 599) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(811 DOWNTO 811)
									);
MUX_REORD_UPDATE_812 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(812 DOWNTO 812) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(601 DOWNTO 601) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(601 DOWNTO 601) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(812 DOWNTO 812)
									);
MUX_REORD_UPDATE_813 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(603 DOWNTO 603) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(603 DOWNTO 603) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(813 DOWNTO 813)
									);
MUX_REORD_UPDATE_814 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(814 DOWNTO 814) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(605 DOWNTO 605) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(605 DOWNTO 605) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(814 DOWNTO 814)
									);
MUX_REORD_UPDATE_815 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(607 DOWNTO 607) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(607 DOWNTO 607) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(815 DOWNTO 815)
									);
MUX_REORD_UPDATE_816 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(816 DOWNTO 816) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(609 DOWNTO 609) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(609 DOWNTO 609) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(816 DOWNTO 816)
									);
MUX_REORD_UPDATE_817 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(611 DOWNTO 611) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(611 DOWNTO 611) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(817 DOWNTO 817)
									);
MUX_REORD_UPDATE_818 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(818 DOWNTO 818) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(613 DOWNTO 613) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(613 DOWNTO 613) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(818 DOWNTO 818)
									);
MUX_REORD_UPDATE_819 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(615 DOWNTO 615) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(615 DOWNTO 615) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(819 DOWNTO 819)
									);
MUX_REORD_UPDATE_820 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(820 DOWNTO 820) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(617 DOWNTO 617) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(617 DOWNTO 617) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(820 DOWNTO 820)
									);
MUX_REORD_UPDATE_821 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(619 DOWNTO 619) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(619 DOWNTO 619) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(821 DOWNTO 821)
									);
MUX_REORD_UPDATE_822 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(822 DOWNTO 822) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(621 DOWNTO 621) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(621 DOWNTO 621) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(822 DOWNTO 822)
									);
MUX_REORD_UPDATE_823 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(623 DOWNTO 623) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(623 DOWNTO 623) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(823 DOWNTO 823)
									);
MUX_REORD_UPDATE_824 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(824 DOWNTO 824) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(625 DOWNTO 625) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(625 DOWNTO 625) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(824 DOWNTO 824)
									);
MUX_REORD_UPDATE_825 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(627 DOWNTO 627) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(627 DOWNTO 627) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(825 DOWNTO 825)
									);
MUX_REORD_UPDATE_826 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(826 DOWNTO 826) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(629 DOWNTO 629) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(629 DOWNTO 629) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(826 DOWNTO 826)
									);
MUX_REORD_UPDATE_827 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(631 DOWNTO 631) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(631 DOWNTO 631) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(827 DOWNTO 827)
									);
MUX_REORD_UPDATE_828 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(828 DOWNTO 828) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(633 DOWNTO 633) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(633 DOWNTO 633) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(828 DOWNTO 828)
									);
MUX_REORD_UPDATE_829 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(635 DOWNTO 635) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(635 DOWNTO 635) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(829 DOWNTO 829)
									);
MUX_REORD_UPDATE_830 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(830 DOWNTO 830) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(637 DOWNTO 637) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(637 DOWNTO 637) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(830 DOWNTO 830)
									);
MUX_REORD_UPDATE_831 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(639 DOWNTO 639) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(639 DOWNTO 639) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(831 DOWNTO 831)
									);
MUX_REORD_UPDATE_832 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(832 DOWNTO 832) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(641 DOWNTO 641) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(641 DOWNTO 641) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(832 DOWNTO 832)
									);
MUX_REORD_UPDATE_833 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(643 DOWNTO 643) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(643 DOWNTO 643) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(833 DOWNTO 833)
									);
MUX_REORD_UPDATE_834 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(834 DOWNTO 834) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(645 DOWNTO 645) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(645 DOWNTO 645) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(834 DOWNTO 834)
									);
MUX_REORD_UPDATE_835 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(647 DOWNTO 647) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(647 DOWNTO 647) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(835 DOWNTO 835)
									);
MUX_REORD_UPDATE_836 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(836 DOWNTO 836) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(649 DOWNTO 649) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(649 DOWNTO 649) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(836 DOWNTO 836)
									);
MUX_REORD_UPDATE_837 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(651 DOWNTO 651) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(651 DOWNTO 651) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(837 DOWNTO 837)
									);
MUX_REORD_UPDATE_838 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(838 DOWNTO 838) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(653 DOWNTO 653) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(653 DOWNTO 653) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(838 DOWNTO 838)
									);
MUX_REORD_UPDATE_839 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(655 DOWNTO 655) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(655 DOWNTO 655) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(839 DOWNTO 839)
									);
MUX_REORD_UPDATE_840 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(840 DOWNTO 840) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(657 DOWNTO 657) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(657 DOWNTO 657) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(840 DOWNTO 840)
									);
MUX_REORD_UPDATE_841 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(659 DOWNTO 659) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(659 DOWNTO 659) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(841 DOWNTO 841)
									);
MUX_REORD_UPDATE_842 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(842 DOWNTO 842) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(661 DOWNTO 661) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(661 DOWNTO 661) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(842 DOWNTO 842)
									);
MUX_REORD_UPDATE_843 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(663 DOWNTO 663) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(663 DOWNTO 663) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(843 DOWNTO 843)
									);
MUX_REORD_UPDATE_844 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(844 DOWNTO 844) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(665 DOWNTO 665) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(665 DOWNTO 665) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(844 DOWNTO 844)
									);
MUX_REORD_UPDATE_845 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(667 DOWNTO 667) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(667 DOWNTO 667) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(845 DOWNTO 845)
									);
MUX_REORD_UPDATE_846 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(846 DOWNTO 846) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(669 DOWNTO 669) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(669 DOWNTO 669) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(846 DOWNTO 846)
									);
MUX_REORD_UPDATE_847 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(671 DOWNTO 671) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(671 DOWNTO 671) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(847 DOWNTO 847)
									);
MUX_REORD_UPDATE_848 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(848 DOWNTO 848) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(673 DOWNTO 673) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(673 DOWNTO 673) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(848 DOWNTO 848)
									);
MUX_REORD_UPDATE_849 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(675 DOWNTO 675) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(675 DOWNTO 675) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(849 DOWNTO 849)
									);
MUX_REORD_UPDATE_850 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(850 DOWNTO 850) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(677 DOWNTO 677) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(677 DOWNTO 677) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(850 DOWNTO 850)
									);
MUX_REORD_UPDATE_851 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(679 DOWNTO 679) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(679 DOWNTO 679) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(851 DOWNTO 851)
									);
MUX_REORD_UPDATE_852 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(852 DOWNTO 852) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(681 DOWNTO 681) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(681 DOWNTO 681) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(852 DOWNTO 852)
									);
MUX_REORD_UPDATE_853 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(683 DOWNTO 683) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(683 DOWNTO 683) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(853 DOWNTO 853)
									);
MUX_REORD_UPDATE_854 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(854 DOWNTO 854) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(685 DOWNTO 685) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(685 DOWNTO 685) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(854 DOWNTO 854)
									);
MUX_REORD_UPDATE_855 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(687 DOWNTO 687) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(687 DOWNTO 687) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(855 DOWNTO 855)
									);
MUX_REORD_UPDATE_856 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(856 DOWNTO 856) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(689 DOWNTO 689) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(689 DOWNTO 689) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(856 DOWNTO 856)
									);
MUX_REORD_UPDATE_857 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(691 DOWNTO 691) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(691 DOWNTO 691) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(857 DOWNTO 857)
									);
MUX_REORD_UPDATE_858 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(858 DOWNTO 858) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(693 DOWNTO 693) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(693 DOWNTO 693) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(858 DOWNTO 858)
									);
MUX_REORD_UPDATE_859 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(695 DOWNTO 695) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(695 DOWNTO 695) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(859 DOWNTO 859)
									);
MUX_REORD_UPDATE_860 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(860 DOWNTO 860) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(697 DOWNTO 697) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(697 DOWNTO 697) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(860 DOWNTO 860)
									);
MUX_REORD_UPDATE_861 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(699 DOWNTO 699) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(699 DOWNTO 699) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(861 DOWNTO 861)
									);
MUX_REORD_UPDATE_862 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(862 DOWNTO 862) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(701 DOWNTO 701) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(701 DOWNTO 701) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(862 DOWNTO 862)
									);
MUX_REORD_UPDATE_863 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(703 DOWNTO 703) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(703 DOWNTO 703) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(863 DOWNTO 863)
									);
MUX_REORD_UPDATE_864 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(864 DOWNTO 864) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(705 DOWNTO 705) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(705 DOWNTO 705) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(864 DOWNTO 864)
									);
MUX_REORD_UPDATE_865 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(707 DOWNTO 707) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(707 DOWNTO 707) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(865 DOWNTO 865)
									);
MUX_REORD_UPDATE_866 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(866 DOWNTO 866) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(709 DOWNTO 709) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(709 DOWNTO 709) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(866 DOWNTO 866)
									);
MUX_REORD_UPDATE_867 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(711 DOWNTO 711) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(711 DOWNTO 711) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(867 DOWNTO 867)
									);
MUX_REORD_UPDATE_868 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(868 DOWNTO 868) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(713 DOWNTO 713) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(713 DOWNTO 713) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(868 DOWNTO 868)
									);
MUX_REORD_UPDATE_869 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(715 DOWNTO 715) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(715 DOWNTO 715) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(869 DOWNTO 869)
									);
MUX_REORD_UPDATE_870 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(870 DOWNTO 870) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(717 DOWNTO 717) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(717 DOWNTO 717) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(870 DOWNTO 870)
									);
MUX_REORD_UPDATE_871 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(719 DOWNTO 719) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(719 DOWNTO 719) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(871 DOWNTO 871)
									);
MUX_REORD_UPDATE_872 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(872 DOWNTO 872) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(721 DOWNTO 721) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(721 DOWNTO 721) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(872 DOWNTO 872)
									);
MUX_REORD_UPDATE_873 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(723 DOWNTO 723) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(723 DOWNTO 723) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(873 DOWNTO 873)
									);
MUX_REORD_UPDATE_874 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(874 DOWNTO 874) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(725 DOWNTO 725) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(725 DOWNTO 725) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(874 DOWNTO 874)
									);
MUX_REORD_UPDATE_875 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(727 DOWNTO 727) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(727 DOWNTO 727) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(875 DOWNTO 875)
									);
MUX_REORD_UPDATE_876 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(876 DOWNTO 876) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(729 DOWNTO 729) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(729 DOWNTO 729) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(876 DOWNTO 876)
									);
MUX_REORD_UPDATE_877 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(731 DOWNTO 731) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(731 DOWNTO 731) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(877 DOWNTO 877)
									);
MUX_REORD_UPDATE_878 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(878 DOWNTO 878) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(733 DOWNTO 733) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(733 DOWNTO 733) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(878 DOWNTO 878)
									);
MUX_REORD_UPDATE_879 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(735 DOWNTO 735) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(735 DOWNTO 735) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(879 DOWNTO 879)
									);
MUX_REORD_UPDATE_880 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(880 DOWNTO 880) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(737 DOWNTO 737) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(737 DOWNTO 737) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(880 DOWNTO 880)
									);
MUX_REORD_UPDATE_881 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(739 DOWNTO 739) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(739 DOWNTO 739) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(881 DOWNTO 881)
									);
MUX_REORD_UPDATE_882 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(882 DOWNTO 882) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(741 DOWNTO 741) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(741 DOWNTO 741) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(882 DOWNTO 882)
									);
MUX_REORD_UPDATE_883 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(743 DOWNTO 743) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(743 DOWNTO 743) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(883 DOWNTO 883)
									);
MUX_REORD_UPDATE_884 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(884 DOWNTO 884) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(745 DOWNTO 745) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(745 DOWNTO 745) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(884 DOWNTO 884)
									);
MUX_REORD_UPDATE_885 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(747 DOWNTO 747) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(747 DOWNTO 747) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(885 DOWNTO 885)
									);
MUX_REORD_UPDATE_886 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(886 DOWNTO 886) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(749 DOWNTO 749) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(749 DOWNTO 749) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(886 DOWNTO 886)
									);
MUX_REORD_UPDATE_887 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(751 DOWNTO 751) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(751 DOWNTO 751) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(887 DOWNTO 887)
									);
MUX_REORD_UPDATE_888 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(888 DOWNTO 888) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(753 DOWNTO 753) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(753 DOWNTO 753) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(888 DOWNTO 888)
									);
MUX_REORD_UPDATE_889 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(755 DOWNTO 755) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(755 DOWNTO 755) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(889 DOWNTO 889)
									);
MUX_REORD_UPDATE_890 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(890 DOWNTO 890) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(757 DOWNTO 757) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(757 DOWNTO 757) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(890 DOWNTO 890)
									);
MUX_REORD_UPDATE_891 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(759 DOWNTO 759) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(759 DOWNTO 759) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(891 DOWNTO 891)
									);
MUX_REORD_UPDATE_892 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(892 DOWNTO 892) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(761 DOWNTO 761) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(761 DOWNTO 761) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(892 DOWNTO 892)
									);
MUX_REORD_UPDATE_893 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(763 DOWNTO 763) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(763 DOWNTO 763) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(893 DOWNTO 893)
									);
MUX_REORD_UPDATE_894 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(894 DOWNTO 894) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(765 DOWNTO 765) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(765 DOWNTO 765) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(894 DOWNTO 894)
									);
MUX_REORD_UPDATE_895 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(767 DOWNTO 767) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(767 DOWNTO 767) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(895 DOWNTO 895)
									);
MUX_REORD_UPDATE_896 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(896 DOWNTO 896) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(769 DOWNTO 769) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(769 DOWNTO 769) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(896 DOWNTO 896)
									);
MUX_REORD_UPDATE_897 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(771 DOWNTO 771) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(771 DOWNTO 771) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(897 DOWNTO 897)
									);
MUX_REORD_UPDATE_898 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(898 DOWNTO 898) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(773 DOWNTO 773) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(773 DOWNTO 773) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(898 DOWNTO 898)
									);
MUX_REORD_UPDATE_899 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(775 DOWNTO 775) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(775 DOWNTO 775) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(899 DOWNTO 899)
									);
MUX_REORD_UPDATE_900 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(900 DOWNTO 900) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(777 DOWNTO 777) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(777 DOWNTO 777) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(900 DOWNTO 900)
									);
MUX_REORD_UPDATE_901 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(779 DOWNTO 779) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(779 DOWNTO 779) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(901 DOWNTO 901)
									);
MUX_REORD_UPDATE_902 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(902 DOWNTO 902) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(781 DOWNTO 781) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(781 DOWNTO 781) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(902 DOWNTO 902)
									);
MUX_REORD_UPDATE_903 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(783 DOWNTO 783) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(783 DOWNTO 783) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(903 DOWNTO 903)
									);
MUX_REORD_UPDATE_904 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(904 DOWNTO 904) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(785 DOWNTO 785) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(785 DOWNTO 785) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(904 DOWNTO 904)
									);
MUX_REORD_UPDATE_905 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(787 DOWNTO 787) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(787 DOWNTO 787) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(905 DOWNTO 905)
									);
MUX_REORD_UPDATE_906 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(906 DOWNTO 906) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(789 DOWNTO 789) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(789 DOWNTO 789) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(906 DOWNTO 906)
									);
MUX_REORD_UPDATE_907 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(791 DOWNTO 791) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(791 DOWNTO 791) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(907 DOWNTO 907)
									);
MUX_REORD_UPDATE_908 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(908 DOWNTO 908) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(793 DOWNTO 793) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(793 DOWNTO 793) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(908 DOWNTO 908)
									);
MUX_REORD_UPDATE_909 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(795 DOWNTO 795) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(795 DOWNTO 795) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(909 DOWNTO 909)
									);
MUX_REORD_UPDATE_910 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(910 DOWNTO 910) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(797 DOWNTO 797) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(797 DOWNTO 797) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(910 DOWNTO 910)
									);
MUX_REORD_UPDATE_911 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(799 DOWNTO 799) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(799 DOWNTO 799) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(911 DOWNTO 911)
									);
MUX_REORD_UPDATE_912 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(912 DOWNTO 912) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(801 DOWNTO 801) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(801 DOWNTO 801) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(912 DOWNTO 912)
									);
MUX_REORD_UPDATE_913 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(803 DOWNTO 803) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(803 DOWNTO 803) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(913 DOWNTO 913)
									);
MUX_REORD_UPDATE_914 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(914 DOWNTO 914) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(805 DOWNTO 805) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(805 DOWNTO 805) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(914 DOWNTO 914)
									);
MUX_REORD_UPDATE_915 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(807 DOWNTO 807) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(807 DOWNTO 807) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(915 DOWNTO 915)
									);
MUX_REORD_UPDATE_916 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(916 DOWNTO 916) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(809 DOWNTO 809) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(809 DOWNTO 809) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(916 DOWNTO 916)
									);
MUX_REORD_UPDATE_917 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(811 DOWNTO 811) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(811 DOWNTO 811) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(917 DOWNTO 917)
									);
MUX_REORD_UPDATE_918 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(918 DOWNTO 918) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(813 DOWNTO 813) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(813 DOWNTO 813) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(918 DOWNTO 918)
									);
MUX_REORD_UPDATE_919 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(815 DOWNTO 815) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(815 DOWNTO 815) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(919 DOWNTO 919)
									);
MUX_REORD_UPDATE_920 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(920 DOWNTO 920) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(817 DOWNTO 817) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(817 DOWNTO 817) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(920 DOWNTO 920)
									);
MUX_REORD_UPDATE_921 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(819 DOWNTO 819) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(819 DOWNTO 819) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(921 DOWNTO 921)
									);
MUX_REORD_UPDATE_922 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(922 DOWNTO 922) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(821 DOWNTO 821) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(821 DOWNTO 821) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(922 DOWNTO 922)
									);
MUX_REORD_UPDATE_923 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(823 DOWNTO 823) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(823 DOWNTO 823) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(923 DOWNTO 923)
									);
MUX_REORD_UPDATE_924 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(924 DOWNTO 924) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(825 DOWNTO 825) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(825 DOWNTO 825) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(924 DOWNTO 924)
									);
MUX_REORD_UPDATE_925 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(827 DOWNTO 827) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(827 DOWNTO 827) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(925 DOWNTO 925)
									);
MUX_REORD_UPDATE_926 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(926 DOWNTO 926) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(829 DOWNTO 829) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(829 DOWNTO 829) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(926 DOWNTO 926)
									);
MUX_REORD_UPDATE_927 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(831 DOWNTO 831) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(831 DOWNTO 831) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(927 DOWNTO 927)
									);
MUX_REORD_UPDATE_928 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(928 DOWNTO 928) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(833 DOWNTO 833) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(833 DOWNTO 833) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(928 DOWNTO 928)
									);
MUX_REORD_UPDATE_929 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(835 DOWNTO 835) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(835 DOWNTO 835) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(929 DOWNTO 929)
									);
MUX_REORD_UPDATE_930 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(930 DOWNTO 930) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(837 DOWNTO 837) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(837 DOWNTO 837) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(930 DOWNTO 930)
									);
MUX_REORD_UPDATE_931 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(839 DOWNTO 839) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(839 DOWNTO 839) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(931 DOWNTO 931)
									);
MUX_REORD_UPDATE_932 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(932 DOWNTO 932) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(841 DOWNTO 841) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(841 DOWNTO 841) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(932 DOWNTO 932)
									);
MUX_REORD_UPDATE_933 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(843 DOWNTO 843) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(843 DOWNTO 843) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(933 DOWNTO 933)
									);
MUX_REORD_UPDATE_934 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(934 DOWNTO 934) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(845 DOWNTO 845) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(845 DOWNTO 845) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(934 DOWNTO 934)
									);
MUX_REORD_UPDATE_935 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(847 DOWNTO 847) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(847 DOWNTO 847) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(935 DOWNTO 935)
									);
MUX_REORD_UPDATE_936 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(936 DOWNTO 936) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(849 DOWNTO 849) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(849 DOWNTO 849) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(936 DOWNTO 936)
									);
MUX_REORD_UPDATE_937 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(851 DOWNTO 851) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(851 DOWNTO 851) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(937 DOWNTO 937)
									);
MUX_REORD_UPDATE_938 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(938 DOWNTO 938) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(853 DOWNTO 853) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(853 DOWNTO 853) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(938 DOWNTO 938)
									);
MUX_REORD_UPDATE_939 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(855 DOWNTO 855) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(855 DOWNTO 855) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(939 DOWNTO 939)
									);
MUX_REORD_UPDATE_940 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(940 DOWNTO 940) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(857 DOWNTO 857) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(857 DOWNTO 857) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(940 DOWNTO 940)
									);
MUX_REORD_UPDATE_941 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(859 DOWNTO 859) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(859 DOWNTO 859) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(941 DOWNTO 941)
									);
MUX_REORD_UPDATE_942 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(942 DOWNTO 942) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(861 DOWNTO 861) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(861 DOWNTO 861) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(942 DOWNTO 942)
									);
MUX_REORD_UPDATE_943 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(863 DOWNTO 863) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(863 DOWNTO 863) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(943 DOWNTO 943)
									);
MUX_REORD_UPDATE_944 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(944 DOWNTO 944) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(865 DOWNTO 865) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(865 DOWNTO 865) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(944 DOWNTO 944)
									);
MUX_REORD_UPDATE_945 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(867 DOWNTO 867) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(867 DOWNTO 867) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(945 DOWNTO 945)
									);
MUX_REORD_UPDATE_946 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(946 DOWNTO 946) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(869 DOWNTO 869) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(869 DOWNTO 869) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(946 DOWNTO 946)
									);
MUX_REORD_UPDATE_947 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(871 DOWNTO 871) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(871 DOWNTO 871) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(947 DOWNTO 947)
									);
MUX_REORD_UPDATE_948 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(948 DOWNTO 948) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(873 DOWNTO 873) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(873 DOWNTO 873) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(948 DOWNTO 948)
									);
MUX_REORD_UPDATE_949 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(875 DOWNTO 875) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(875 DOWNTO 875) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(949 DOWNTO 949)
									);
MUX_REORD_UPDATE_950 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(950 DOWNTO 950) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(877 DOWNTO 877) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(877 DOWNTO 877) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(950 DOWNTO 950)
									);
MUX_REORD_UPDATE_951 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(879 DOWNTO 879) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(879 DOWNTO 879) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(951 DOWNTO 951)
									);
MUX_REORD_UPDATE_952 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(952 DOWNTO 952) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(881 DOWNTO 881) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(881 DOWNTO 881) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(952 DOWNTO 952)
									);
MUX_REORD_UPDATE_953 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(883 DOWNTO 883) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(883 DOWNTO 883) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(953 DOWNTO 953)
									);
MUX_REORD_UPDATE_954 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(954 DOWNTO 954) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(885 DOWNTO 885) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(885 DOWNTO 885) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(954 DOWNTO 954)
									);
MUX_REORD_UPDATE_955 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(887 DOWNTO 887) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(887 DOWNTO 887) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(955 DOWNTO 955)
									);
MUX_REORD_UPDATE_956 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(956 DOWNTO 956) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(889 DOWNTO 889) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(889 DOWNTO 889) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(956 DOWNTO 956)
									);
MUX_REORD_UPDATE_957 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(891 DOWNTO 891) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(891 DOWNTO 891) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(957 DOWNTO 957)
									);
MUX_REORD_UPDATE_958 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(958 DOWNTO 958) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(893 DOWNTO 893) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(893 DOWNTO 893) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(958 DOWNTO 958)
									);
MUX_REORD_UPDATE_959 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(895 DOWNTO 895) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(895 DOWNTO 895) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(959 DOWNTO 959)
									);
MUX_REORD_UPDATE_960 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(960 DOWNTO 960) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(897 DOWNTO 897) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(897 DOWNTO 897) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(960 DOWNTO 960)
									);
MUX_REORD_UPDATE_961 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(899 DOWNTO 899) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(899 DOWNTO 899) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(961 DOWNTO 961)
									);
MUX_REORD_UPDATE_962 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(962 DOWNTO 962) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(901 DOWNTO 901) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(901 DOWNTO 901) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(962 DOWNTO 962)
									);
MUX_REORD_UPDATE_963 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(903 DOWNTO 903) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(903 DOWNTO 903) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(963 DOWNTO 963)
									);
MUX_REORD_UPDATE_964 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(964 DOWNTO 964) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(905 DOWNTO 905) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(905 DOWNTO 905) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(964 DOWNTO 964)
									);
MUX_REORD_UPDATE_965 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(907 DOWNTO 907) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(907 DOWNTO 907) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(965 DOWNTO 965)
									);
MUX_REORD_UPDATE_966 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(966 DOWNTO 966) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(909 DOWNTO 909) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(909 DOWNTO 909) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(966 DOWNTO 966)
									);
MUX_REORD_UPDATE_967 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(911 DOWNTO 911) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(911 DOWNTO 911) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(967 DOWNTO 967)
									);
MUX_REORD_UPDATE_968 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(968 DOWNTO 968) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(913 DOWNTO 913) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(913 DOWNTO 913) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(968 DOWNTO 968)
									);
MUX_REORD_UPDATE_969 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(915 DOWNTO 915) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(915 DOWNTO 915) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(969 DOWNTO 969)
									);
MUX_REORD_UPDATE_970 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(970 DOWNTO 970) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(917 DOWNTO 917) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(917 DOWNTO 917) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(970 DOWNTO 970)
									);
MUX_REORD_UPDATE_971 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(919 DOWNTO 919) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(919 DOWNTO 919) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(971 DOWNTO 971)
									);
MUX_REORD_UPDATE_972 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(972 DOWNTO 972) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(921 DOWNTO 921) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(921 DOWNTO 921) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(972 DOWNTO 972)
									);
MUX_REORD_UPDATE_973 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(923 DOWNTO 923) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(923 DOWNTO 923) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(973 DOWNTO 973)
									);
MUX_REORD_UPDATE_974 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(974 DOWNTO 974) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(925 DOWNTO 925) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(925 DOWNTO 925) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(974 DOWNTO 974)
									);
MUX_REORD_UPDATE_975 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(927 DOWNTO 927) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(927 DOWNTO 927) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(975 DOWNTO 975)
									);
MUX_REORD_UPDATE_976 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(976 DOWNTO 976) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(929 DOWNTO 929) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(929 DOWNTO 929) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(976 DOWNTO 976)
									);
MUX_REORD_UPDATE_977 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(931 DOWNTO 931) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(931 DOWNTO 931) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(977 DOWNTO 977)
									);
MUX_REORD_UPDATE_978 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(978 DOWNTO 978) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(933 DOWNTO 933) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(933 DOWNTO 933) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(978 DOWNTO 978)
									);
MUX_REORD_UPDATE_979 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(935 DOWNTO 935) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(935 DOWNTO 935) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(979 DOWNTO 979)
									);
MUX_REORD_UPDATE_980 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(980 DOWNTO 980) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(937 DOWNTO 937) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(937 DOWNTO 937) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(980 DOWNTO 980)
									);
MUX_REORD_UPDATE_981 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(939 DOWNTO 939) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(939 DOWNTO 939) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(981 DOWNTO 981)
									);
MUX_REORD_UPDATE_982 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(982 DOWNTO 982) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(941 DOWNTO 941) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(941 DOWNTO 941) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(982 DOWNTO 982)
									);
MUX_REORD_UPDATE_983 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(943 DOWNTO 943) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(943 DOWNTO 943) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(983 DOWNTO 983)
									);
MUX_REORD_UPDATE_984 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(984 DOWNTO 984) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(945 DOWNTO 945) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(945 DOWNTO 945) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(984 DOWNTO 984)
									);
MUX_REORD_UPDATE_985 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(947 DOWNTO 947) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(947 DOWNTO 947) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(985 DOWNTO 985)
									);
MUX_REORD_UPDATE_986 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(986 DOWNTO 986) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(949 DOWNTO 949) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(949 DOWNTO 949) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(986 DOWNTO 986)
									);
MUX_REORD_UPDATE_987 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(951 DOWNTO 951) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(951 DOWNTO 951) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(987 DOWNTO 987)
									);
MUX_REORD_UPDATE_988 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(988 DOWNTO 988) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(953 DOWNTO 953) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(953 DOWNTO 953) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(988 DOWNTO 988)
									);
MUX_REORD_UPDATE_989 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(955 DOWNTO 955) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(955 DOWNTO 955) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(989 DOWNTO 989)
									);
MUX_REORD_UPDATE_990 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(990 DOWNTO 990) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(957 DOWNTO 957) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(957 DOWNTO 957) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(990 DOWNTO 990)
									);
MUX_REORD_UPDATE_991 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(959 DOWNTO 959) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(959 DOWNTO 959) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(991 DOWNTO 991)
									);
MUX_REORD_UPDATE_992 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(992 DOWNTO 992) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(961 DOWNTO 961) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(961 DOWNTO 961) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(992 DOWNTO 992)
									);
MUX_REORD_UPDATE_993 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(963 DOWNTO 963) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(963 DOWNTO 963) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(993 DOWNTO 993)
									);
MUX_REORD_UPDATE_994 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(994 DOWNTO 994) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(965 DOWNTO 965) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(965 DOWNTO 965) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(994 DOWNTO 994)
									);
MUX_REORD_UPDATE_995 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(967 DOWNTO 967) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(967 DOWNTO 967) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(995 DOWNTO 995)
									);
MUX_REORD_UPDATE_996 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(996 DOWNTO 996) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(969 DOWNTO 969) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(969 DOWNTO 969) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(996 DOWNTO 996)
									);
MUX_REORD_UPDATE_997 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(971 DOWNTO 971) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(971 DOWNTO 971) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(997 DOWNTO 997)
									);
MUX_REORD_UPDATE_998 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(998 DOWNTO 998) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(973 DOWNTO 973) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(973 DOWNTO 973) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(998 DOWNTO 998)
									);
MUX_REORD_UPDATE_999 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(975 DOWNTO 975) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(975 DOWNTO 975) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(999 DOWNTO 999)
									);
MUX_REORD_UPDATE_1000 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1000 DOWNTO 1000) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(977 DOWNTO 977) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(977 DOWNTO 977) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1000 DOWNTO 1000)
									);
MUX_REORD_UPDATE_1001 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(979 DOWNTO 979) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(979 DOWNTO 979) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1001 DOWNTO 1001)
									);
MUX_REORD_UPDATE_1002 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1002 DOWNTO 1002) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(981 DOWNTO 981) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(981 DOWNTO 981) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1002 DOWNTO 1002)
									);
MUX_REORD_UPDATE_1003 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(983 DOWNTO 983) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(983 DOWNTO 983) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1003 DOWNTO 1003)
									);
MUX_REORD_UPDATE_1004 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1004 DOWNTO 1004) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(985 DOWNTO 985) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(985 DOWNTO 985) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1004 DOWNTO 1004)
									);
MUX_REORD_UPDATE_1005 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(987 DOWNTO 987) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(987 DOWNTO 987) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1005 DOWNTO 1005)
									);
MUX_REORD_UPDATE_1006 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1006 DOWNTO 1006) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(989 DOWNTO 989) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(989 DOWNTO 989) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1006 DOWNTO 1006)
									);
MUX_REORD_UPDATE_1007 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(991 DOWNTO 991) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(991 DOWNTO 991) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1007 DOWNTO 1007)
									);
MUX_REORD_UPDATE_1008 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1008 DOWNTO 1008) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(993 DOWNTO 993) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(993 DOWNTO 993) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1008 DOWNTO 1008)
									);
MUX_REORD_UPDATE_1009 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(995 DOWNTO 995) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(995 DOWNTO 995) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1009 DOWNTO 1009)
									);
MUX_REORD_UPDATE_1010 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1010 DOWNTO 1010) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(997 DOWNTO 997) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(997 DOWNTO 997) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1010 DOWNTO 1010)
									);
MUX_REORD_UPDATE_1011 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(999 DOWNTO 999) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(999 DOWNTO 999) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1011 DOWNTO 1011)
									);
MUX_REORD_UPDATE_1012 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1012 DOWNTO 1012) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1001 DOWNTO 1001) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1012 DOWNTO 1012)
									);
MUX_REORD_UPDATE_1013 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1003 DOWNTO 1003) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1013 DOWNTO 1013)
									);
MUX_REORD_UPDATE_1014 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1014 DOWNTO 1014) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1005 DOWNTO 1005) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1014 DOWNTO 1014)
									);
MUX_REORD_UPDATE_1015 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1007 DOWNTO 1007) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1015 DOWNTO 1015)
									);
MUX_REORD_UPDATE_1016 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1016 DOWNTO 1016) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1009 DOWNTO 1009) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1016 DOWNTO 1016)
									);
MUX_REORD_UPDATE_1017 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1011 DOWNTO 1011) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1017 DOWNTO 1017)
									);
MUX_REORD_UPDATE_1018 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1018 DOWNTO 1018) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1013 DOWNTO 1013) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1018 DOWNTO 1018)
									);
MUX_REORD_UPDATE_1019 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1015 DOWNTO 1015) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1019 DOWNTO 1019)
									);
MUX_REORD_UPDATE_1020 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1020 DOWNTO 1020) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1017 DOWNTO 1017) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1020 DOWNTO 1020)
									);
MUX_REORD_UPDATE_1021 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1019 DOWNTO 1019) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1021 DOWNTO 1021)
									);
MUX_REORD_UPDATE_1022 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1022 DOWNTO 1022) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1021 DOWNTO 1021) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1022 DOWNTO 1022)
									);
MUX_REORD_UPDATE_1023 : multiplexer_10_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_1 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_2 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_3 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_4 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_5 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_6 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_7 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_8 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
										MUX_10_1_IN_9 => UNWINDOWED_MASK(1023 DOWNTO 1023) ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => REORDERED_MASK(1023 DOWNTO 1023)
									);

STATE_UPDATE_MASK(0) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(0) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(0);
STATE_UPDATE_MASK(1) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1);
STATE_UPDATE_MASK(2) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(2) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(2);
STATE_UPDATE_MASK(3) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(3) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(3);
STATE_UPDATE_MASK(4) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(4) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(4);
STATE_UPDATE_MASK(5) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(5) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(5);
STATE_UPDATE_MASK(6) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(6) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(6);
STATE_UPDATE_MASK(7) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(7) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(7);
STATE_UPDATE_MASK(8) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(8) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(8);
STATE_UPDATE_MASK(9) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(9) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(9);
STATE_UPDATE_MASK(10) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(10) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(10);
STATE_UPDATE_MASK(11) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(11) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(11);
STATE_UPDATE_MASK(12) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(12) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(12);
STATE_UPDATE_MASK(13) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(13) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(13);
STATE_UPDATE_MASK(14) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(14) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(14);
STATE_UPDATE_MASK(15) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(15) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(15);
STATE_UPDATE_MASK(16) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(16) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(16);
STATE_UPDATE_MASK(17) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(17) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(17);
STATE_UPDATE_MASK(18) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(18) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(18);
STATE_UPDATE_MASK(19) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(19) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(19);
STATE_UPDATE_MASK(20) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(20) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(20);
STATE_UPDATE_MASK(21) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(21) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(21);
STATE_UPDATE_MASK(22) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(22) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(22);
STATE_UPDATE_MASK(23) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(23) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(23);
STATE_UPDATE_MASK(24) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(24) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(24);
STATE_UPDATE_MASK(25) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(25) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(25);
STATE_UPDATE_MASK(26) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(26) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(26);
STATE_UPDATE_MASK(27) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(27) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(27);
STATE_UPDATE_MASK(28) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(28) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(28);
STATE_UPDATE_MASK(29) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(29) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(29);
STATE_UPDATE_MASK(30) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(30) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(30);
STATE_UPDATE_MASK(31) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(31) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(31);
STATE_UPDATE_MASK(32) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(32) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(32);
STATE_UPDATE_MASK(33) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(33) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(33);
STATE_UPDATE_MASK(34) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(34) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(34);
STATE_UPDATE_MASK(35) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(35) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(35);
STATE_UPDATE_MASK(36) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(36) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(36);
STATE_UPDATE_MASK(37) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(37) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(37);
STATE_UPDATE_MASK(38) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(38) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(38);
STATE_UPDATE_MASK(39) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(39) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(39);
STATE_UPDATE_MASK(40) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(40) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(40);
STATE_UPDATE_MASK(41) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(41) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(41);
STATE_UPDATE_MASK(42) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(42) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(42);
STATE_UPDATE_MASK(43) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(43) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(43);
STATE_UPDATE_MASK(44) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(44) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(44);
STATE_UPDATE_MASK(45) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(45) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(45);
STATE_UPDATE_MASK(46) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(46) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(46);
STATE_UPDATE_MASK(47) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(47) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(47);
STATE_UPDATE_MASK(48) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(48) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(48);
STATE_UPDATE_MASK(49) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(49) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(49);
STATE_UPDATE_MASK(50) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(50) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(50);
STATE_UPDATE_MASK(51) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(51) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(51);
STATE_UPDATE_MASK(52) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(52) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(52);
STATE_UPDATE_MASK(53) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(53) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(53);
STATE_UPDATE_MASK(54) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(54) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(54);
STATE_UPDATE_MASK(55) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(55) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(55);
STATE_UPDATE_MASK(56) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(56) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(56);
STATE_UPDATE_MASK(57) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(57) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(57);
STATE_UPDATE_MASK(58) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(58) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(58);
STATE_UPDATE_MASK(59) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(59) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(59);
STATE_UPDATE_MASK(60) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(60) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(60);
STATE_UPDATE_MASK(61) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(61) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(61);
STATE_UPDATE_MASK(62) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(62) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(62);
STATE_UPDATE_MASK(63) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(63) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(63);
STATE_UPDATE_MASK(64) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(64) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(64);
STATE_UPDATE_MASK(65) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(65) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(65);
STATE_UPDATE_MASK(66) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(66) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(66);
STATE_UPDATE_MASK(67) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(67) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(67);
STATE_UPDATE_MASK(68) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(68) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(68);
STATE_UPDATE_MASK(69) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(69) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(69);
STATE_UPDATE_MASK(70) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(70) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(70);
STATE_UPDATE_MASK(71) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(71) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(71);
STATE_UPDATE_MASK(72) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(72) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(72);
STATE_UPDATE_MASK(73) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(73) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(73);
STATE_UPDATE_MASK(74) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(74) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(74);
STATE_UPDATE_MASK(75) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(75) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(75);
STATE_UPDATE_MASK(76) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(76) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(76);
STATE_UPDATE_MASK(77) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(77) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(77);
STATE_UPDATE_MASK(78) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(78) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(78);
STATE_UPDATE_MASK(79) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(79) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(79);
STATE_UPDATE_MASK(80) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(80) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(80);
STATE_UPDATE_MASK(81) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(81) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(81);
STATE_UPDATE_MASK(82) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(82) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(82);
STATE_UPDATE_MASK(83) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(83) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(83);
STATE_UPDATE_MASK(84) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(84) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(84);
STATE_UPDATE_MASK(85) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(85) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(85);
STATE_UPDATE_MASK(86) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(86) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(86);
STATE_UPDATE_MASK(87) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(87) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(87);
STATE_UPDATE_MASK(88) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(88) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(88);
STATE_UPDATE_MASK(89) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(89) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(89);
STATE_UPDATE_MASK(90) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(90) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(90);
STATE_UPDATE_MASK(91) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(91) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(91);
STATE_UPDATE_MASK(92) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(92) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(92);
STATE_UPDATE_MASK(93) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(93) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(93);
STATE_UPDATE_MASK(94) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(94) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(94);
STATE_UPDATE_MASK(95) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(95) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(95);
STATE_UPDATE_MASK(96) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(96) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(96);
STATE_UPDATE_MASK(97) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(97) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(97);
STATE_UPDATE_MASK(98) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(98) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(98);
STATE_UPDATE_MASK(99) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(99) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(99);
STATE_UPDATE_MASK(100) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(100) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(100);
STATE_UPDATE_MASK(101) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(101) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(101);
STATE_UPDATE_MASK(102) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(102) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(102);
STATE_UPDATE_MASK(103) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(103) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(103);
STATE_UPDATE_MASK(104) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(104) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(104);
STATE_UPDATE_MASK(105) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(105) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(105);
STATE_UPDATE_MASK(106) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(106) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(106);
STATE_UPDATE_MASK(107) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(107) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(107);
STATE_UPDATE_MASK(108) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(108) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(108);
STATE_UPDATE_MASK(109) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(109) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(109);
STATE_UPDATE_MASK(110) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(110) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(110);
STATE_UPDATE_MASK(111) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(111) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(111);
STATE_UPDATE_MASK(112) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(112) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(112);
STATE_UPDATE_MASK(113) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(113) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(113);
STATE_UPDATE_MASK(114) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(114) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(114);
STATE_UPDATE_MASK(115) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(115) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(115);
STATE_UPDATE_MASK(116) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(116) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(116);
STATE_UPDATE_MASK(117) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(117) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(117);
STATE_UPDATE_MASK(118) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(118) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(118);
STATE_UPDATE_MASK(119) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(119) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(119);
STATE_UPDATE_MASK(120) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(120) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(120);
STATE_UPDATE_MASK(121) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(121) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(121);
STATE_UPDATE_MASK(122) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(122) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(122);
STATE_UPDATE_MASK(123) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(123) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(123);
STATE_UPDATE_MASK(124) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(124) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(124);
STATE_UPDATE_MASK(125) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(125) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(125);
STATE_UPDATE_MASK(126) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(126) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(126);
STATE_UPDATE_MASK(127) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(127) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(127);
STATE_UPDATE_MASK(128) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(128) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(128);
STATE_UPDATE_MASK(129) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(129) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(129);
STATE_UPDATE_MASK(130) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(130) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(130);
STATE_UPDATE_MASK(131) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(131) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(131);
STATE_UPDATE_MASK(132) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(132) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(132);
STATE_UPDATE_MASK(133) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(133) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(133);
STATE_UPDATE_MASK(134) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(134) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(134);
STATE_UPDATE_MASK(135) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(135) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(135);
STATE_UPDATE_MASK(136) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(136) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(136);
STATE_UPDATE_MASK(137) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(137) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(137);
STATE_UPDATE_MASK(138) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(138) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(138);
STATE_UPDATE_MASK(139) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(139) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(139);
STATE_UPDATE_MASK(140) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(140) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(140);
STATE_UPDATE_MASK(141) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(141) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(141);
STATE_UPDATE_MASK(142) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(142) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(142);
STATE_UPDATE_MASK(143) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(143) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(143);
STATE_UPDATE_MASK(144) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(144) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(144);
STATE_UPDATE_MASK(145) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(145) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(145);
STATE_UPDATE_MASK(146) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(146) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(146);
STATE_UPDATE_MASK(147) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(147) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(147);
STATE_UPDATE_MASK(148) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(148) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(148);
STATE_UPDATE_MASK(149) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(149) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(149);
STATE_UPDATE_MASK(150) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(150) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(150);
STATE_UPDATE_MASK(151) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(151) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(151);
STATE_UPDATE_MASK(152) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(152) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(152);
STATE_UPDATE_MASK(153) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(153) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(153);
STATE_UPDATE_MASK(154) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(154) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(154);
STATE_UPDATE_MASK(155) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(155) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(155);
STATE_UPDATE_MASK(156) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(156) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(156);
STATE_UPDATE_MASK(157) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(157) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(157);
STATE_UPDATE_MASK(158) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(158) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(158);
STATE_UPDATE_MASK(159) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(159) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(159);
STATE_UPDATE_MASK(160) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(160) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(160);
STATE_UPDATE_MASK(161) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(161) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(161);
STATE_UPDATE_MASK(162) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(162) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(162);
STATE_UPDATE_MASK(163) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(163) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(163);
STATE_UPDATE_MASK(164) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(164) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(164);
STATE_UPDATE_MASK(165) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(165) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(165);
STATE_UPDATE_MASK(166) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(166) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(166);
STATE_UPDATE_MASK(167) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(167) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(167);
STATE_UPDATE_MASK(168) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(168) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(168);
STATE_UPDATE_MASK(169) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(169) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(169);
STATE_UPDATE_MASK(170) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(170) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(170);
STATE_UPDATE_MASK(171) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(171) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(171);
STATE_UPDATE_MASK(172) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(172) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(172);
STATE_UPDATE_MASK(173) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(173) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(173);
STATE_UPDATE_MASK(174) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(174) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(174);
STATE_UPDATE_MASK(175) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(175) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(175);
STATE_UPDATE_MASK(176) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(176) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(176);
STATE_UPDATE_MASK(177) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(177) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(177);
STATE_UPDATE_MASK(178) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(178) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(178);
STATE_UPDATE_MASK(179) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(179) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(179);
STATE_UPDATE_MASK(180) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(180) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(180);
STATE_UPDATE_MASK(181) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(181) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(181);
STATE_UPDATE_MASK(182) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(182) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(182);
STATE_UPDATE_MASK(183) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(183) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(183);
STATE_UPDATE_MASK(184) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(184) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(184);
STATE_UPDATE_MASK(185) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(185) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(185);
STATE_UPDATE_MASK(186) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(186) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(186);
STATE_UPDATE_MASK(187) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(187) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(187);
STATE_UPDATE_MASK(188) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(188) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(188);
STATE_UPDATE_MASK(189) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(189) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(189);
STATE_UPDATE_MASK(190) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(190) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(190);
STATE_UPDATE_MASK(191) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(191) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(191);
STATE_UPDATE_MASK(192) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(192) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(192);
STATE_UPDATE_MASK(193) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(193) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(193);
STATE_UPDATE_MASK(194) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(194) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(194);
STATE_UPDATE_MASK(195) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(195) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(195);
STATE_UPDATE_MASK(196) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(196) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(196);
STATE_UPDATE_MASK(197) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(197) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(197);
STATE_UPDATE_MASK(198) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(198) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(198);
STATE_UPDATE_MASK(199) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(199) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(199);
STATE_UPDATE_MASK(200) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(200) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(200);
STATE_UPDATE_MASK(201) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(201) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(201);
STATE_UPDATE_MASK(202) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(202) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(202);
STATE_UPDATE_MASK(203) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(203) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(203);
STATE_UPDATE_MASK(204) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(204) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(204);
STATE_UPDATE_MASK(205) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(205) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(205);
STATE_UPDATE_MASK(206) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(206) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(206);
STATE_UPDATE_MASK(207) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(207) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(207);
STATE_UPDATE_MASK(208) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(208) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(208);
STATE_UPDATE_MASK(209) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(209) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(209);
STATE_UPDATE_MASK(210) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(210) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(210);
STATE_UPDATE_MASK(211) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(211) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(211);
STATE_UPDATE_MASK(212) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(212) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(212);
STATE_UPDATE_MASK(213) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(213) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(213);
STATE_UPDATE_MASK(214) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(214) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(214);
STATE_UPDATE_MASK(215) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(215) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(215);
STATE_UPDATE_MASK(216) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(216) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(216);
STATE_UPDATE_MASK(217) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(217) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(217);
STATE_UPDATE_MASK(218) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(218) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(218);
STATE_UPDATE_MASK(219) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(219) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(219);
STATE_UPDATE_MASK(220) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(220) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(220);
STATE_UPDATE_MASK(221) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(221) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(221);
STATE_UPDATE_MASK(222) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(222) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(222);
STATE_UPDATE_MASK(223) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(223) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(223);
STATE_UPDATE_MASK(224) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(224) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(224);
STATE_UPDATE_MASK(225) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(225) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(225);
STATE_UPDATE_MASK(226) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(226) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(226);
STATE_UPDATE_MASK(227) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(227) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(227);
STATE_UPDATE_MASK(228) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(228) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(228);
STATE_UPDATE_MASK(229) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(229) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(229);
STATE_UPDATE_MASK(230) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(230) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(230);
STATE_UPDATE_MASK(231) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(231) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(231);
STATE_UPDATE_MASK(232) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(232) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(232);
STATE_UPDATE_MASK(233) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(233) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(233);
STATE_UPDATE_MASK(234) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(234) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(234);
STATE_UPDATE_MASK(235) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(235) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(235);
STATE_UPDATE_MASK(236) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(236) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(236);
STATE_UPDATE_MASK(237) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(237) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(237);
STATE_UPDATE_MASK(238) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(238) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(238);
STATE_UPDATE_MASK(239) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(239) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(239);
STATE_UPDATE_MASK(240) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(240) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(240);
STATE_UPDATE_MASK(241) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(241) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(241);
STATE_UPDATE_MASK(242) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(242) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(242);
STATE_UPDATE_MASK(243) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(243) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(243);
STATE_UPDATE_MASK(244) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(244) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(244);
STATE_UPDATE_MASK(245) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(245) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(245);
STATE_UPDATE_MASK(246) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(246) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(246);
STATE_UPDATE_MASK(247) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(247) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(247);
STATE_UPDATE_MASK(248) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(248) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(248);
STATE_UPDATE_MASK(249) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(249) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(249);
STATE_UPDATE_MASK(250) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(250) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(250);
STATE_UPDATE_MASK(251) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(251) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(251);
STATE_UPDATE_MASK(252) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(252) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(252);
STATE_UPDATE_MASK(253) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(253) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(253);
STATE_UPDATE_MASK(254) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(254) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(254);
STATE_UPDATE_MASK(255) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(255) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(255);
STATE_UPDATE_MASK(256) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(256) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(256);
STATE_UPDATE_MASK(257) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(257) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(257);
STATE_UPDATE_MASK(258) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(258) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(258);
STATE_UPDATE_MASK(259) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(259) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(259);
STATE_UPDATE_MASK(260) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(260) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(260);
STATE_UPDATE_MASK(261) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(261) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(261);
STATE_UPDATE_MASK(262) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(262) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(262);
STATE_UPDATE_MASK(263) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(263) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(263);
STATE_UPDATE_MASK(264) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(264) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(264);
STATE_UPDATE_MASK(265) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(265) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(265);
STATE_UPDATE_MASK(266) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(266) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(266);
STATE_UPDATE_MASK(267) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(267) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(267);
STATE_UPDATE_MASK(268) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(268) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(268);
STATE_UPDATE_MASK(269) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(269) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(269);
STATE_UPDATE_MASK(270) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(270) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(270);
STATE_UPDATE_MASK(271) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(271) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(271);
STATE_UPDATE_MASK(272) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(272) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(272);
STATE_UPDATE_MASK(273) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(273) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(273);
STATE_UPDATE_MASK(274) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(274) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(274);
STATE_UPDATE_MASK(275) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(275) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(275);
STATE_UPDATE_MASK(276) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(276) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(276);
STATE_UPDATE_MASK(277) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(277) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(277);
STATE_UPDATE_MASK(278) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(278) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(278);
STATE_UPDATE_MASK(279) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(279) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(279);
STATE_UPDATE_MASK(280) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(280) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(280);
STATE_UPDATE_MASK(281) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(281) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(281);
STATE_UPDATE_MASK(282) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(282) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(282);
STATE_UPDATE_MASK(283) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(283) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(283);
STATE_UPDATE_MASK(284) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(284) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(284);
STATE_UPDATE_MASK(285) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(285) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(285);
STATE_UPDATE_MASK(286) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(286) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(286);
STATE_UPDATE_MASK(287) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(287) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(287);
STATE_UPDATE_MASK(288) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(288) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(288);
STATE_UPDATE_MASK(289) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(289) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(289);
STATE_UPDATE_MASK(290) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(290) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(290);
STATE_UPDATE_MASK(291) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(291) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(291);
STATE_UPDATE_MASK(292) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(292) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(292);
STATE_UPDATE_MASK(293) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(293) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(293);
STATE_UPDATE_MASK(294) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(294) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(294);
STATE_UPDATE_MASK(295) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(295) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(295);
STATE_UPDATE_MASK(296) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(296) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(296);
STATE_UPDATE_MASK(297) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(297) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(297);
STATE_UPDATE_MASK(298) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(298) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(298);
STATE_UPDATE_MASK(299) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(299) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(299);
STATE_UPDATE_MASK(300) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(300) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(300);
STATE_UPDATE_MASK(301) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(301) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(301);
STATE_UPDATE_MASK(302) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(302) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(302);
STATE_UPDATE_MASK(303) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(303) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(303);
STATE_UPDATE_MASK(304) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(304) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(304);
STATE_UPDATE_MASK(305) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(305) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(305);
STATE_UPDATE_MASK(306) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(306) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(306);
STATE_UPDATE_MASK(307) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(307) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(307);
STATE_UPDATE_MASK(308) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(308) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(308);
STATE_UPDATE_MASK(309) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(309) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(309);
STATE_UPDATE_MASK(310) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(310) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(310);
STATE_UPDATE_MASK(311) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(311) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(311);
STATE_UPDATE_MASK(312) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(312) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(312);
STATE_UPDATE_MASK(313) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(313) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(313);
STATE_UPDATE_MASK(314) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(314) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(314);
STATE_UPDATE_MASK(315) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(315) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(315);
STATE_UPDATE_MASK(316) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(316) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(316);
STATE_UPDATE_MASK(317) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(317) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(317);
STATE_UPDATE_MASK(318) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(318) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(318);
STATE_UPDATE_MASK(319) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(319) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(319);
STATE_UPDATE_MASK(320) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(320) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(320);
STATE_UPDATE_MASK(321) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(321) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(321);
STATE_UPDATE_MASK(322) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(322) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(322);
STATE_UPDATE_MASK(323) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(323) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(323);
STATE_UPDATE_MASK(324) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(324) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(324);
STATE_UPDATE_MASK(325) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(325) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(325);
STATE_UPDATE_MASK(326) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(326) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(326);
STATE_UPDATE_MASK(327) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(327) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(327);
STATE_UPDATE_MASK(328) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(328) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(328);
STATE_UPDATE_MASK(329) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(329) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(329);
STATE_UPDATE_MASK(330) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(330) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(330);
STATE_UPDATE_MASK(331) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(331) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(331);
STATE_UPDATE_MASK(332) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(332) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(332);
STATE_UPDATE_MASK(333) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(333) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(333);
STATE_UPDATE_MASK(334) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(334) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(334);
STATE_UPDATE_MASK(335) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(335) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(335);
STATE_UPDATE_MASK(336) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(336) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(336);
STATE_UPDATE_MASK(337) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(337) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(337);
STATE_UPDATE_MASK(338) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(338) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(338);
STATE_UPDATE_MASK(339) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(339) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(339);
STATE_UPDATE_MASK(340) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(340) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(340);
STATE_UPDATE_MASK(341) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(341) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(341);
STATE_UPDATE_MASK(342) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(342) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(342);
STATE_UPDATE_MASK(343) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(343) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(343);
STATE_UPDATE_MASK(344) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(344) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(344);
STATE_UPDATE_MASK(345) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(345) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(345);
STATE_UPDATE_MASK(346) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(346) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(346);
STATE_UPDATE_MASK(347) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(347) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(347);
STATE_UPDATE_MASK(348) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(348) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(348);
STATE_UPDATE_MASK(349) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(349) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(349);
STATE_UPDATE_MASK(350) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(350) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(350);
STATE_UPDATE_MASK(351) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(351) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(351);
STATE_UPDATE_MASK(352) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(352) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(352);
STATE_UPDATE_MASK(353) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(353) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(353);
STATE_UPDATE_MASK(354) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(354) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(354);
STATE_UPDATE_MASK(355) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(355) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(355);
STATE_UPDATE_MASK(356) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(356) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(356);
STATE_UPDATE_MASK(357) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(357) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(357);
STATE_UPDATE_MASK(358) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(358) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(358);
STATE_UPDATE_MASK(359) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(359) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(359);
STATE_UPDATE_MASK(360) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(360) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(360);
STATE_UPDATE_MASK(361) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(361) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(361);
STATE_UPDATE_MASK(362) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(362) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(362);
STATE_UPDATE_MASK(363) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(363) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(363);
STATE_UPDATE_MASK(364) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(364) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(364);
STATE_UPDATE_MASK(365) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(365) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(365);
STATE_UPDATE_MASK(366) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(366) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(366);
STATE_UPDATE_MASK(367) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(367) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(367);
STATE_UPDATE_MASK(368) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(368) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(368);
STATE_UPDATE_MASK(369) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(369) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(369);
STATE_UPDATE_MASK(370) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(370) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(370);
STATE_UPDATE_MASK(371) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(371) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(371);
STATE_UPDATE_MASK(372) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(372) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(372);
STATE_UPDATE_MASK(373) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(373) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(373);
STATE_UPDATE_MASK(374) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(374) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(374);
STATE_UPDATE_MASK(375) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(375) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(375);
STATE_UPDATE_MASK(376) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(376) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(376);
STATE_UPDATE_MASK(377) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(377) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(377);
STATE_UPDATE_MASK(378) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(378) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(378);
STATE_UPDATE_MASK(379) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(379) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(379);
STATE_UPDATE_MASK(380) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(380) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(380);
STATE_UPDATE_MASK(381) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(381) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(381);
STATE_UPDATE_MASK(382) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(382) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(382);
STATE_UPDATE_MASK(383) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(383) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(383);
STATE_UPDATE_MASK(384) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(384) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(384);
STATE_UPDATE_MASK(385) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(385) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(385);
STATE_UPDATE_MASK(386) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(386) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(386);
STATE_UPDATE_MASK(387) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(387) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(387);
STATE_UPDATE_MASK(388) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(388) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(388);
STATE_UPDATE_MASK(389) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(389) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(389);
STATE_UPDATE_MASK(390) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(390) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(390);
STATE_UPDATE_MASK(391) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(391) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(391);
STATE_UPDATE_MASK(392) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(392) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(392);
STATE_UPDATE_MASK(393) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(393) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(393);
STATE_UPDATE_MASK(394) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(394) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(394);
STATE_UPDATE_MASK(395) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(395) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(395);
STATE_UPDATE_MASK(396) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(396) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(396);
STATE_UPDATE_MASK(397) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(397) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(397);
STATE_UPDATE_MASK(398) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(398) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(398);
STATE_UPDATE_MASK(399) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(399) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(399);
STATE_UPDATE_MASK(400) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(400) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(400);
STATE_UPDATE_MASK(401) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(401) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(401);
STATE_UPDATE_MASK(402) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(402) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(402);
STATE_UPDATE_MASK(403) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(403) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(403);
STATE_UPDATE_MASK(404) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(404) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(404);
STATE_UPDATE_MASK(405) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(405) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(405);
STATE_UPDATE_MASK(406) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(406) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(406);
STATE_UPDATE_MASK(407) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(407) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(407);
STATE_UPDATE_MASK(408) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(408) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(408);
STATE_UPDATE_MASK(409) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(409) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(409);
STATE_UPDATE_MASK(410) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(410) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(410);
STATE_UPDATE_MASK(411) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(411) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(411);
STATE_UPDATE_MASK(412) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(412) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(412);
STATE_UPDATE_MASK(413) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(413) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(413);
STATE_UPDATE_MASK(414) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(414) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(414);
STATE_UPDATE_MASK(415) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(415) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(415);
STATE_UPDATE_MASK(416) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(416) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(416);
STATE_UPDATE_MASK(417) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(417) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(417);
STATE_UPDATE_MASK(418) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(418) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(418);
STATE_UPDATE_MASK(419) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(419) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(419);
STATE_UPDATE_MASK(420) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(420) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(420);
STATE_UPDATE_MASK(421) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(421) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(421);
STATE_UPDATE_MASK(422) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(422) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(422);
STATE_UPDATE_MASK(423) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(423) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(423);
STATE_UPDATE_MASK(424) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(424) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(424);
STATE_UPDATE_MASK(425) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(425) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(425);
STATE_UPDATE_MASK(426) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(426) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(426);
STATE_UPDATE_MASK(427) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(427) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(427);
STATE_UPDATE_MASK(428) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(428) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(428);
STATE_UPDATE_MASK(429) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(429) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(429);
STATE_UPDATE_MASK(430) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(430) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(430);
STATE_UPDATE_MASK(431) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(431) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(431);
STATE_UPDATE_MASK(432) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(432) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(432);
STATE_UPDATE_MASK(433) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(433) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(433);
STATE_UPDATE_MASK(434) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(434) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(434);
STATE_UPDATE_MASK(435) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(435) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(435);
STATE_UPDATE_MASK(436) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(436) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(436);
STATE_UPDATE_MASK(437) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(437) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(437);
STATE_UPDATE_MASK(438) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(438) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(438);
STATE_UPDATE_MASK(439) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(439) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(439);
STATE_UPDATE_MASK(440) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(440) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(440);
STATE_UPDATE_MASK(441) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(441) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(441);
STATE_UPDATE_MASK(442) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(442) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(442);
STATE_UPDATE_MASK(443) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(443) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(443);
STATE_UPDATE_MASK(444) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(444) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(444);
STATE_UPDATE_MASK(445) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(445) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(445);
STATE_UPDATE_MASK(446) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(446) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(446);
STATE_UPDATE_MASK(447) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(447) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(447);
STATE_UPDATE_MASK(448) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(448) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(448);
STATE_UPDATE_MASK(449) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(449) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(449);
STATE_UPDATE_MASK(450) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(450) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(450);
STATE_UPDATE_MASK(451) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(451) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(451);
STATE_UPDATE_MASK(452) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(452) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(452);
STATE_UPDATE_MASK(453) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(453) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(453);
STATE_UPDATE_MASK(454) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(454) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(454);
STATE_UPDATE_MASK(455) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(455) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(455);
STATE_UPDATE_MASK(456) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(456) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(456);
STATE_UPDATE_MASK(457) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(457) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(457);
STATE_UPDATE_MASK(458) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(458) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(458);
STATE_UPDATE_MASK(459) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(459) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(459);
STATE_UPDATE_MASK(460) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(460) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(460);
STATE_UPDATE_MASK(461) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(461) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(461);
STATE_UPDATE_MASK(462) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(462) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(462);
STATE_UPDATE_MASK(463) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(463) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(463);
STATE_UPDATE_MASK(464) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(464) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(464);
STATE_UPDATE_MASK(465) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(465) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(465);
STATE_UPDATE_MASK(466) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(466) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(466);
STATE_UPDATE_MASK(467) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(467) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(467);
STATE_UPDATE_MASK(468) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(468) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(468);
STATE_UPDATE_MASK(469) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(469) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(469);
STATE_UPDATE_MASK(470) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(470) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(470);
STATE_UPDATE_MASK(471) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(471) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(471);
STATE_UPDATE_MASK(472) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(472) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(472);
STATE_UPDATE_MASK(473) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(473) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(473);
STATE_UPDATE_MASK(474) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(474) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(474);
STATE_UPDATE_MASK(475) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(475) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(475);
STATE_UPDATE_MASK(476) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(476) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(476);
STATE_UPDATE_MASK(477) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(477) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(477);
STATE_UPDATE_MASK(478) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(478) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(478);
STATE_UPDATE_MASK(479) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(479) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(479);
STATE_UPDATE_MASK(480) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(480) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(480);
STATE_UPDATE_MASK(481) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(481) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(481);
STATE_UPDATE_MASK(482) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(482) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(482);
STATE_UPDATE_MASK(483) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(483) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(483);
STATE_UPDATE_MASK(484) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(484) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(484);
STATE_UPDATE_MASK(485) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(485) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(485);
STATE_UPDATE_MASK(486) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(486) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(486);
STATE_UPDATE_MASK(487) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(487) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(487);
STATE_UPDATE_MASK(488) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(488) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(488);
STATE_UPDATE_MASK(489) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(489) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(489);
STATE_UPDATE_MASK(490) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(490) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(490);
STATE_UPDATE_MASK(491) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(491) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(491);
STATE_UPDATE_MASK(492) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(492) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(492);
STATE_UPDATE_MASK(493) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(493) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(493);
STATE_UPDATE_MASK(494) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(494) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(494);
STATE_UPDATE_MASK(495) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(495) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(495);
STATE_UPDATE_MASK(496) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(496) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(496);
STATE_UPDATE_MASK(497) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(497) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(497);
STATE_UPDATE_MASK(498) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(498) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(498);
STATE_UPDATE_MASK(499) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(499) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(499);
STATE_UPDATE_MASK(500) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(500) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(500);
STATE_UPDATE_MASK(501) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(501) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(501);
STATE_UPDATE_MASK(502) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(502) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(502);
STATE_UPDATE_MASK(503) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(503) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(503);
STATE_UPDATE_MASK(504) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(504) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(504);
STATE_UPDATE_MASK(505) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(505) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(505);
STATE_UPDATE_MASK(506) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(506) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(506);
STATE_UPDATE_MASK(507) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(507) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(507);
STATE_UPDATE_MASK(508) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(508) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(508);
STATE_UPDATE_MASK(509) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(509) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(509);
STATE_UPDATE_MASK(510) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(510) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(510);
STATE_UPDATE_MASK(511) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(511) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(511);
STATE_UPDATE_MASK(512) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(512) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(512);
STATE_UPDATE_MASK(513) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(513) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(513);
STATE_UPDATE_MASK(514) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(514) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(514);
STATE_UPDATE_MASK(515) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(515) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(515);
STATE_UPDATE_MASK(516) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(516) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(516);
STATE_UPDATE_MASK(517) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(517) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(517);
STATE_UPDATE_MASK(518) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(518) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(518);
STATE_UPDATE_MASK(519) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(519) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(519);
STATE_UPDATE_MASK(520) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(520) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(520);
STATE_UPDATE_MASK(521) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(521) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(521);
STATE_UPDATE_MASK(522) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(522) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(522);
STATE_UPDATE_MASK(523) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(523) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(523);
STATE_UPDATE_MASK(524) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(524) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(524);
STATE_UPDATE_MASK(525) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(525) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(525);
STATE_UPDATE_MASK(526) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(526) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(526);
STATE_UPDATE_MASK(527) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(527) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(527);
STATE_UPDATE_MASK(528) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(528) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(528);
STATE_UPDATE_MASK(529) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(529) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(529);
STATE_UPDATE_MASK(530) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(530) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(530);
STATE_UPDATE_MASK(531) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(531) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(531);
STATE_UPDATE_MASK(532) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(532) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(532);
STATE_UPDATE_MASK(533) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(533) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(533);
STATE_UPDATE_MASK(534) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(534) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(534);
STATE_UPDATE_MASK(535) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(535) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(535);
STATE_UPDATE_MASK(536) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(536) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(536);
STATE_UPDATE_MASK(537) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(537) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(537);
STATE_UPDATE_MASK(538) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(538) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(538);
STATE_UPDATE_MASK(539) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(539) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(539);
STATE_UPDATE_MASK(540) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(540) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(540);
STATE_UPDATE_MASK(541) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(541) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(541);
STATE_UPDATE_MASK(542) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(542) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(542);
STATE_UPDATE_MASK(543) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(543) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(543);
STATE_UPDATE_MASK(544) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(544) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(544);
STATE_UPDATE_MASK(545) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(545) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(545);
STATE_UPDATE_MASK(546) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(546) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(546);
STATE_UPDATE_MASK(547) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(547) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(547);
STATE_UPDATE_MASK(548) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(548) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(548);
STATE_UPDATE_MASK(549) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(549) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(549);
STATE_UPDATE_MASK(550) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(550) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(550);
STATE_UPDATE_MASK(551) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(551) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(551);
STATE_UPDATE_MASK(552) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(552) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(552);
STATE_UPDATE_MASK(553) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(553) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(553);
STATE_UPDATE_MASK(554) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(554) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(554);
STATE_UPDATE_MASK(555) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(555) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(555);
STATE_UPDATE_MASK(556) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(556) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(556);
STATE_UPDATE_MASK(557) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(557) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(557);
STATE_UPDATE_MASK(558) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(558) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(558);
STATE_UPDATE_MASK(559) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(559) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(559);
STATE_UPDATE_MASK(560) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(560) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(560);
STATE_UPDATE_MASK(561) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(561) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(561);
STATE_UPDATE_MASK(562) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(562) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(562);
STATE_UPDATE_MASK(563) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(563) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(563);
STATE_UPDATE_MASK(564) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(564) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(564);
STATE_UPDATE_MASK(565) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(565) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(565);
STATE_UPDATE_MASK(566) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(566) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(566);
STATE_UPDATE_MASK(567) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(567) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(567);
STATE_UPDATE_MASK(568) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(568) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(568);
STATE_UPDATE_MASK(569) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(569) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(569);
STATE_UPDATE_MASK(570) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(570) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(570);
STATE_UPDATE_MASK(571) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(571) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(571);
STATE_UPDATE_MASK(572) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(572) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(572);
STATE_UPDATE_MASK(573) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(573) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(573);
STATE_UPDATE_MASK(574) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(574) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(574);
STATE_UPDATE_MASK(575) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(575) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(575);
STATE_UPDATE_MASK(576) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(576) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(576);
STATE_UPDATE_MASK(577) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(577) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(577);
STATE_UPDATE_MASK(578) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(578) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(578);
STATE_UPDATE_MASK(579) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(579) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(579);
STATE_UPDATE_MASK(580) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(580) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(580);
STATE_UPDATE_MASK(581) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(581) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(581);
STATE_UPDATE_MASK(582) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(582) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(582);
STATE_UPDATE_MASK(583) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(583) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(583);
STATE_UPDATE_MASK(584) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(584) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(584);
STATE_UPDATE_MASK(585) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(585) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(585);
STATE_UPDATE_MASK(586) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(586) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(586);
STATE_UPDATE_MASK(587) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(587) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(587);
STATE_UPDATE_MASK(588) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(588) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(588);
STATE_UPDATE_MASK(589) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(589) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(589);
STATE_UPDATE_MASK(590) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(590) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(590);
STATE_UPDATE_MASK(591) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(591) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(591);
STATE_UPDATE_MASK(592) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(592) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(592);
STATE_UPDATE_MASK(593) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(593) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(593);
STATE_UPDATE_MASK(594) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(594) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(594);
STATE_UPDATE_MASK(595) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(595) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(595);
STATE_UPDATE_MASK(596) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(596) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(596);
STATE_UPDATE_MASK(597) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(597) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(597);
STATE_UPDATE_MASK(598) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(598) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(598);
STATE_UPDATE_MASK(599) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(599) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(599);
STATE_UPDATE_MASK(600) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(600) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(600);
STATE_UPDATE_MASK(601) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(601) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(601);
STATE_UPDATE_MASK(602) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(602) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(602);
STATE_UPDATE_MASK(603) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(603) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(603);
STATE_UPDATE_MASK(604) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(604) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(604);
STATE_UPDATE_MASK(605) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(605) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(605);
STATE_UPDATE_MASK(606) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(606) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(606);
STATE_UPDATE_MASK(607) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(607) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(607);
STATE_UPDATE_MASK(608) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(608) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(608);
STATE_UPDATE_MASK(609) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(609) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(609);
STATE_UPDATE_MASK(610) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(610) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(610);
STATE_UPDATE_MASK(611) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(611) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(611);
STATE_UPDATE_MASK(612) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(612) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(612);
STATE_UPDATE_MASK(613) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(613) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(613);
STATE_UPDATE_MASK(614) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(614) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(614);
STATE_UPDATE_MASK(615) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(615) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(615);
STATE_UPDATE_MASK(616) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(616) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(616);
STATE_UPDATE_MASK(617) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(617) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(617);
STATE_UPDATE_MASK(618) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(618) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(618);
STATE_UPDATE_MASK(619) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(619) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(619);
STATE_UPDATE_MASK(620) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(620) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(620);
STATE_UPDATE_MASK(621) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(621) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(621);
STATE_UPDATE_MASK(622) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(622) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(622);
STATE_UPDATE_MASK(623) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(623) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(623);
STATE_UPDATE_MASK(624) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(624) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(624);
STATE_UPDATE_MASK(625) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(625) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(625);
STATE_UPDATE_MASK(626) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(626) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(626);
STATE_UPDATE_MASK(627) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(627) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(627);
STATE_UPDATE_MASK(628) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(628) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(628);
STATE_UPDATE_MASK(629) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(629) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(629);
STATE_UPDATE_MASK(630) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(630) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(630);
STATE_UPDATE_MASK(631) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(631) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(631);
STATE_UPDATE_MASK(632) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(632) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(632);
STATE_UPDATE_MASK(633) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(633) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(633);
STATE_UPDATE_MASK(634) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(634) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(634);
STATE_UPDATE_MASK(635) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(635) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(635);
STATE_UPDATE_MASK(636) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(636) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(636);
STATE_UPDATE_MASK(637) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(637) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(637);
STATE_UPDATE_MASK(638) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(638) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(638);
STATE_UPDATE_MASK(639) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(639) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(639);
STATE_UPDATE_MASK(640) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(640) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(640);
STATE_UPDATE_MASK(641) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(641) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(641);
STATE_UPDATE_MASK(642) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(642) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(642);
STATE_UPDATE_MASK(643) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(643) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(643);
STATE_UPDATE_MASK(644) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(644) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(644);
STATE_UPDATE_MASK(645) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(645) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(645);
STATE_UPDATE_MASK(646) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(646) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(646);
STATE_UPDATE_MASK(647) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(647) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(647);
STATE_UPDATE_MASK(648) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(648) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(648);
STATE_UPDATE_MASK(649) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(649) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(649);
STATE_UPDATE_MASK(650) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(650) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(650);
STATE_UPDATE_MASK(651) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(651) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(651);
STATE_UPDATE_MASK(652) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(652) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(652);
STATE_UPDATE_MASK(653) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(653) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(653);
STATE_UPDATE_MASK(654) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(654) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(654);
STATE_UPDATE_MASK(655) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(655) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(655);
STATE_UPDATE_MASK(656) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(656) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(656);
STATE_UPDATE_MASK(657) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(657) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(657);
STATE_UPDATE_MASK(658) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(658) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(658);
STATE_UPDATE_MASK(659) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(659) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(659);
STATE_UPDATE_MASK(660) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(660) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(660);
STATE_UPDATE_MASK(661) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(661) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(661);
STATE_UPDATE_MASK(662) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(662) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(662);
STATE_UPDATE_MASK(663) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(663) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(663);
STATE_UPDATE_MASK(664) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(664) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(664);
STATE_UPDATE_MASK(665) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(665) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(665);
STATE_UPDATE_MASK(666) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(666) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(666);
STATE_UPDATE_MASK(667) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(667) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(667);
STATE_UPDATE_MASK(668) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(668) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(668);
STATE_UPDATE_MASK(669) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(669) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(669);
STATE_UPDATE_MASK(670) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(670) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(670);
STATE_UPDATE_MASK(671) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(671) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(671);
STATE_UPDATE_MASK(672) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(672) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(672);
STATE_UPDATE_MASK(673) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(673) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(673);
STATE_UPDATE_MASK(674) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(674) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(674);
STATE_UPDATE_MASK(675) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(675) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(675);
STATE_UPDATE_MASK(676) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(676) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(676);
STATE_UPDATE_MASK(677) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(677) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(677);
STATE_UPDATE_MASK(678) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(678) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(678);
STATE_UPDATE_MASK(679) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(679) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(679);
STATE_UPDATE_MASK(680) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(680) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(680);
STATE_UPDATE_MASK(681) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(681) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(681);
STATE_UPDATE_MASK(682) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(682) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(682);
STATE_UPDATE_MASK(683) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(683) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(683);
STATE_UPDATE_MASK(684) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(684) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(684);
STATE_UPDATE_MASK(685) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(685) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(685);
STATE_UPDATE_MASK(686) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(686) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(686);
STATE_UPDATE_MASK(687) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(687) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(687);
STATE_UPDATE_MASK(688) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(688) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(688);
STATE_UPDATE_MASK(689) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(689) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(689);
STATE_UPDATE_MASK(690) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(690) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(690);
STATE_UPDATE_MASK(691) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(691) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(691);
STATE_UPDATE_MASK(692) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(692) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(692);
STATE_UPDATE_MASK(693) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(693) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(693);
STATE_UPDATE_MASK(694) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(694) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(694);
STATE_UPDATE_MASK(695) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(695) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(695);
STATE_UPDATE_MASK(696) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(696) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(696);
STATE_UPDATE_MASK(697) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(697) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(697);
STATE_UPDATE_MASK(698) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(698) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(698);
STATE_UPDATE_MASK(699) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(699) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(699);
STATE_UPDATE_MASK(700) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(700) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(700);
STATE_UPDATE_MASK(701) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(701) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(701);
STATE_UPDATE_MASK(702) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(702) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(702);
STATE_UPDATE_MASK(703) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(703) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(703);
STATE_UPDATE_MASK(704) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(704) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(704);
STATE_UPDATE_MASK(705) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(705) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(705);
STATE_UPDATE_MASK(706) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(706) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(706);
STATE_UPDATE_MASK(707) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(707) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(707);
STATE_UPDATE_MASK(708) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(708) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(708);
STATE_UPDATE_MASK(709) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(709) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(709);
STATE_UPDATE_MASK(710) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(710) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(710);
STATE_UPDATE_MASK(711) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(711) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(711);
STATE_UPDATE_MASK(712) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(712) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(712);
STATE_UPDATE_MASK(713) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(713) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(713);
STATE_UPDATE_MASK(714) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(714) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(714);
STATE_UPDATE_MASK(715) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(715) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(715);
STATE_UPDATE_MASK(716) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(716) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(716);
STATE_UPDATE_MASK(717) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(717) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(717);
STATE_UPDATE_MASK(718) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(718) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(718);
STATE_UPDATE_MASK(719) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(719) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(719);
STATE_UPDATE_MASK(720) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(720) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(720);
STATE_UPDATE_MASK(721) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(721) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(721);
STATE_UPDATE_MASK(722) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(722) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(722);
STATE_UPDATE_MASK(723) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(723) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(723);
STATE_UPDATE_MASK(724) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(724) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(724);
STATE_UPDATE_MASK(725) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(725) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(725);
STATE_UPDATE_MASK(726) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(726) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(726);
STATE_UPDATE_MASK(727) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(727) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(727);
STATE_UPDATE_MASK(728) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(728) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(728);
STATE_UPDATE_MASK(729) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(729) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(729);
STATE_UPDATE_MASK(730) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(730) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(730);
STATE_UPDATE_MASK(731) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(731) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(731);
STATE_UPDATE_MASK(732) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(732) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(732);
STATE_UPDATE_MASK(733) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(733) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(733);
STATE_UPDATE_MASK(734) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(734) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(734);
STATE_UPDATE_MASK(735) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(735) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(735);
STATE_UPDATE_MASK(736) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(736) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(736);
STATE_UPDATE_MASK(737) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(737) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(737);
STATE_UPDATE_MASK(738) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(738) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(738);
STATE_UPDATE_MASK(739) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(739) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(739);
STATE_UPDATE_MASK(740) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(740) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(740);
STATE_UPDATE_MASK(741) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(741) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(741);
STATE_UPDATE_MASK(742) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(742) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(742);
STATE_UPDATE_MASK(743) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(743) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(743);
STATE_UPDATE_MASK(744) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(744) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(744);
STATE_UPDATE_MASK(745) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(745) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(745);
STATE_UPDATE_MASK(746) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(746) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(746);
STATE_UPDATE_MASK(747) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(747) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(747);
STATE_UPDATE_MASK(748) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(748) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(748);
STATE_UPDATE_MASK(749) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(749) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(749);
STATE_UPDATE_MASK(750) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(750) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(750);
STATE_UPDATE_MASK(751) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(751) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(751);
STATE_UPDATE_MASK(752) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(752) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(752);
STATE_UPDATE_MASK(753) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(753) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(753);
STATE_UPDATE_MASK(754) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(754) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(754);
STATE_UPDATE_MASK(755) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(755) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(755);
STATE_UPDATE_MASK(756) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(756) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(756);
STATE_UPDATE_MASK(757) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(757) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(757);
STATE_UPDATE_MASK(758) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(758) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(758);
STATE_UPDATE_MASK(759) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(759) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(759);
STATE_UPDATE_MASK(760) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(760) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(760);
STATE_UPDATE_MASK(761) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(761) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(761);
STATE_UPDATE_MASK(762) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(762) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(762);
STATE_UPDATE_MASK(763) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(763) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(763);
STATE_UPDATE_MASK(764) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(764) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(764);
STATE_UPDATE_MASK(765) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(765) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(765);
STATE_UPDATE_MASK(766) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(766) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(766);
STATE_UPDATE_MASK(767) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(767) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(767);
STATE_UPDATE_MASK(768) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(768) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(768);
STATE_UPDATE_MASK(769) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(769) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(769);
STATE_UPDATE_MASK(770) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(770) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(770);
STATE_UPDATE_MASK(771) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(771) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(771);
STATE_UPDATE_MASK(772) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(772) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(772);
STATE_UPDATE_MASK(773) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(773) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(773);
STATE_UPDATE_MASK(774) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(774) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(774);
STATE_UPDATE_MASK(775) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(775) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(775);
STATE_UPDATE_MASK(776) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(776) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(776);
STATE_UPDATE_MASK(777) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(777) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(777);
STATE_UPDATE_MASK(778) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(778) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(778);
STATE_UPDATE_MASK(779) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(779) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(779);
STATE_UPDATE_MASK(780) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(780) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(780);
STATE_UPDATE_MASK(781) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(781) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(781);
STATE_UPDATE_MASK(782) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(782) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(782);
STATE_UPDATE_MASK(783) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(783) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(783);
STATE_UPDATE_MASK(784) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(784) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(784);
STATE_UPDATE_MASK(785) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(785) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(785);
STATE_UPDATE_MASK(786) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(786) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(786);
STATE_UPDATE_MASK(787) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(787) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(787);
STATE_UPDATE_MASK(788) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(788) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(788);
STATE_UPDATE_MASK(789) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(789) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(789);
STATE_UPDATE_MASK(790) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(790) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(790);
STATE_UPDATE_MASK(791) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(791) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(791);
STATE_UPDATE_MASK(792) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(792) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(792);
STATE_UPDATE_MASK(793) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(793) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(793);
STATE_UPDATE_MASK(794) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(794) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(794);
STATE_UPDATE_MASK(795) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(795) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(795);
STATE_UPDATE_MASK(796) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(796) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(796);
STATE_UPDATE_MASK(797) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(797) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(797);
STATE_UPDATE_MASK(798) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(798) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(798);
STATE_UPDATE_MASK(799) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(799) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(799);
STATE_UPDATE_MASK(800) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(800) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(800);
STATE_UPDATE_MASK(801) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(801) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(801);
STATE_UPDATE_MASK(802) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(802) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(802);
STATE_UPDATE_MASK(803) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(803) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(803);
STATE_UPDATE_MASK(804) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(804) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(804);
STATE_UPDATE_MASK(805) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(805) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(805);
STATE_UPDATE_MASK(806) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(806) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(806);
STATE_UPDATE_MASK(807) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(807) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(807);
STATE_UPDATE_MASK(808) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(808) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(808);
STATE_UPDATE_MASK(809) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(809) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(809);
STATE_UPDATE_MASK(810) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(810) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(810);
STATE_UPDATE_MASK(811) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(811) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(811);
STATE_UPDATE_MASK(812) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(812) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(812);
STATE_UPDATE_MASK(813) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(813) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(813);
STATE_UPDATE_MASK(814) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(814) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(814);
STATE_UPDATE_MASK(815) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(815) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(815);
STATE_UPDATE_MASK(816) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(816) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(816);
STATE_UPDATE_MASK(817) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(817) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(817);
STATE_UPDATE_MASK(818) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(818) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(818);
STATE_UPDATE_MASK(819) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(819) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(819);
STATE_UPDATE_MASK(820) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(820) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(820);
STATE_UPDATE_MASK(821) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(821) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(821);
STATE_UPDATE_MASK(822) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(822) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(822);
STATE_UPDATE_MASK(823) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(823) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(823);
STATE_UPDATE_MASK(824) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(824) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(824);
STATE_UPDATE_MASK(825) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(825) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(825);
STATE_UPDATE_MASK(826) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(826) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(826);
STATE_UPDATE_MASK(827) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(827) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(827);
STATE_UPDATE_MASK(828) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(828) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(828);
STATE_UPDATE_MASK(829) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(829) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(829);
STATE_UPDATE_MASK(830) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(830) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(830);
STATE_UPDATE_MASK(831) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(831) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(831);
STATE_UPDATE_MASK(832) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(832) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(832);
STATE_UPDATE_MASK(833) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(833) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(833);
STATE_UPDATE_MASK(834) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(834) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(834);
STATE_UPDATE_MASK(835) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(835) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(835);
STATE_UPDATE_MASK(836) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(836) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(836);
STATE_UPDATE_MASK(837) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(837) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(837);
STATE_UPDATE_MASK(838) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(838) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(838);
STATE_UPDATE_MASK(839) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(839) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(839);
STATE_UPDATE_MASK(840) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(840) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(840);
STATE_UPDATE_MASK(841) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(841) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(841);
STATE_UPDATE_MASK(842) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(842) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(842);
STATE_UPDATE_MASK(843) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(843) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(843);
STATE_UPDATE_MASK(844) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(844) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(844);
STATE_UPDATE_MASK(845) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(845) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(845);
STATE_UPDATE_MASK(846) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(846) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(846);
STATE_UPDATE_MASK(847) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(847) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(847);
STATE_UPDATE_MASK(848) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(848) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(848);
STATE_UPDATE_MASK(849) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(849) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(849);
STATE_UPDATE_MASK(850) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(850) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(850);
STATE_UPDATE_MASK(851) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(851) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(851);
STATE_UPDATE_MASK(852) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(852) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(852);
STATE_UPDATE_MASK(853) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(853) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(853);
STATE_UPDATE_MASK(854) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(854) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(854);
STATE_UPDATE_MASK(855) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(855) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(855);
STATE_UPDATE_MASK(856) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(856) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(856);
STATE_UPDATE_MASK(857) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(857) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(857);
STATE_UPDATE_MASK(858) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(858) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(858);
STATE_UPDATE_MASK(859) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(859) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(859);
STATE_UPDATE_MASK(860) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(860) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(860);
STATE_UPDATE_MASK(861) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(861) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(861);
STATE_UPDATE_MASK(862) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(862) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(862);
STATE_UPDATE_MASK(863) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(863) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(863);
STATE_UPDATE_MASK(864) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(864) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(864);
STATE_UPDATE_MASK(865) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(865) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(865);
STATE_UPDATE_MASK(866) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(866) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(866);
STATE_UPDATE_MASK(867) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(867) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(867);
STATE_UPDATE_MASK(868) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(868) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(868);
STATE_UPDATE_MASK(869) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(869) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(869);
STATE_UPDATE_MASK(870) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(870) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(870);
STATE_UPDATE_MASK(871) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(871) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(871);
STATE_UPDATE_MASK(872) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(872) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(872);
STATE_UPDATE_MASK(873) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(873) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(873);
STATE_UPDATE_MASK(874) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(874) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(874);
STATE_UPDATE_MASK(875) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(875) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(875);
STATE_UPDATE_MASK(876) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(876) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(876);
STATE_UPDATE_MASK(877) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(877) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(877);
STATE_UPDATE_MASK(878) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(878) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(878);
STATE_UPDATE_MASK(879) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(879) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(879);
STATE_UPDATE_MASK(880) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(880) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(880);
STATE_UPDATE_MASK(881) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(881) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(881);
STATE_UPDATE_MASK(882) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(882) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(882);
STATE_UPDATE_MASK(883) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(883) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(883);
STATE_UPDATE_MASK(884) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(884) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(884);
STATE_UPDATE_MASK(885) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(885) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(885);
STATE_UPDATE_MASK(886) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(886) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(886);
STATE_UPDATE_MASK(887) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(887) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(887);
STATE_UPDATE_MASK(888) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(888) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(888);
STATE_UPDATE_MASK(889) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(889) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(889);
STATE_UPDATE_MASK(890) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(890) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(890);
STATE_UPDATE_MASK(891) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(891) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(891);
STATE_UPDATE_MASK(892) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(892) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(892);
STATE_UPDATE_MASK(893) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(893) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(893);
STATE_UPDATE_MASK(894) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(894) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(894);
STATE_UPDATE_MASK(895) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(895) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(895);
STATE_UPDATE_MASK(896) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(896) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(896);
STATE_UPDATE_MASK(897) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(897) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(897);
STATE_UPDATE_MASK(898) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(898) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(898);
STATE_UPDATE_MASK(899) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(899) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(899);
STATE_UPDATE_MASK(900) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(900) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(900);
STATE_UPDATE_MASK(901) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(901) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(901);
STATE_UPDATE_MASK(902) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(902) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(902);
STATE_UPDATE_MASK(903) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(903) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(903);
STATE_UPDATE_MASK(904) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(904) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(904);
STATE_UPDATE_MASK(905) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(905) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(905);
STATE_UPDATE_MASK(906) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(906) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(906);
STATE_UPDATE_MASK(907) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(907) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(907);
STATE_UPDATE_MASK(908) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(908) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(908);
STATE_UPDATE_MASK(909) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(909) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(909);
STATE_UPDATE_MASK(910) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(910) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(910);
STATE_UPDATE_MASK(911) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(911) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(911);
STATE_UPDATE_MASK(912) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(912) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(912);
STATE_UPDATE_MASK(913) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(913) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(913);
STATE_UPDATE_MASK(914) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(914) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(914);
STATE_UPDATE_MASK(915) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(915) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(915);
STATE_UPDATE_MASK(916) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(916) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(916);
STATE_UPDATE_MASK(917) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(917) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(917);
STATE_UPDATE_MASK(918) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(918) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(918);
STATE_UPDATE_MASK(919) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(919) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(919);
STATE_UPDATE_MASK(920) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(920) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(920);
STATE_UPDATE_MASK(921) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(921) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(921);
STATE_UPDATE_MASK(922) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(922) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(922);
STATE_UPDATE_MASK(923) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(923) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(923);
STATE_UPDATE_MASK(924) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(924) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(924);
STATE_UPDATE_MASK(925) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(925) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(925);
STATE_UPDATE_MASK(926) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(926) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(926);
STATE_UPDATE_MASK(927) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(927) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(927);
STATE_UPDATE_MASK(928) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(928) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(928);
STATE_UPDATE_MASK(929) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(929) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(929);
STATE_UPDATE_MASK(930) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(930) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(930);
STATE_UPDATE_MASK(931) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(931) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(931);
STATE_UPDATE_MASK(932) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(932) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(932);
STATE_UPDATE_MASK(933) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(933) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(933);
STATE_UPDATE_MASK(934) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(934) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(934);
STATE_UPDATE_MASK(935) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(935) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(935);
STATE_UPDATE_MASK(936) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(936) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(936);
STATE_UPDATE_MASK(937) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(937) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(937);
STATE_UPDATE_MASK(938) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(938) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(938);
STATE_UPDATE_MASK(939) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(939) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(939);
STATE_UPDATE_MASK(940) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(940) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(940);
STATE_UPDATE_MASK(941) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(941) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(941);
STATE_UPDATE_MASK(942) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(942) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(942);
STATE_UPDATE_MASK(943) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(943) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(943);
STATE_UPDATE_MASK(944) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(944) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(944);
STATE_UPDATE_MASK(945) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(945) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(945);
STATE_UPDATE_MASK(946) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(946) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(946);
STATE_UPDATE_MASK(947) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(947) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(947);
STATE_UPDATE_MASK(948) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(948) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(948);
STATE_UPDATE_MASK(949) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(949) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(949);
STATE_UPDATE_MASK(950) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(950) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(950);
STATE_UPDATE_MASK(951) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(951) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(951);
STATE_UPDATE_MASK(952) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(952) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(952);
STATE_UPDATE_MASK(953) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(953) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(953);
STATE_UPDATE_MASK(954) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(954) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(954);
STATE_UPDATE_MASK(955) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(955) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(955);
STATE_UPDATE_MASK(956) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(956) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(956);
STATE_UPDATE_MASK(957) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(957) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(957);
STATE_UPDATE_MASK(958) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(958) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(958);
STATE_UPDATE_MASK(959) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(959) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(959);
STATE_UPDATE_MASK(960) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(960) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(960);
STATE_UPDATE_MASK(961) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(961) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(961);
STATE_UPDATE_MASK(962) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(962) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(962);
STATE_UPDATE_MASK(963) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(963) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(963);
STATE_UPDATE_MASK(964) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(964) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(964);
STATE_UPDATE_MASK(965) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(965) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(965);
STATE_UPDATE_MASK(966) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(966) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(966);
STATE_UPDATE_MASK(967) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(967) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(967);
STATE_UPDATE_MASK(968) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(968) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(968);
STATE_UPDATE_MASK(969) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(969) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(969);
STATE_UPDATE_MASK(970) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(970) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(970);
STATE_UPDATE_MASK(971) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(971) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(971);
STATE_UPDATE_MASK(972) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(972) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(972);
STATE_UPDATE_MASK(973) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(973) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(973);
STATE_UPDATE_MASK(974) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(974) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(974);
STATE_UPDATE_MASK(975) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(975) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(975);
STATE_UPDATE_MASK(976) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(976) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(976);
STATE_UPDATE_MASK(977) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(977) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(977);
STATE_UPDATE_MASK(978) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(978) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(978);
STATE_UPDATE_MASK(979) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(979) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(979);
STATE_UPDATE_MASK(980) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(980) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(980);
STATE_UPDATE_MASK(981) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(981) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(981);
STATE_UPDATE_MASK(982) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(982) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(982);
STATE_UPDATE_MASK(983) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(983) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(983);
STATE_UPDATE_MASK(984) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(984) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(984);
STATE_UPDATE_MASK(985) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(985) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(985);
STATE_UPDATE_MASK(986) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(986) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(986);
STATE_UPDATE_MASK(987) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(987) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(987);
STATE_UPDATE_MASK(988) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(988) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(988);
STATE_UPDATE_MASK(989) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(989) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(989);
STATE_UPDATE_MASK(990) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(990) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(990);
STATE_UPDATE_MASK(991) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(991) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(991);
STATE_UPDATE_MASK(992) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(992) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(992);
STATE_UPDATE_MASK(993) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(993) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(993);
STATE_UPDATE_MASK(994) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(994) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(994);
STATE_UPDATE_MASK(995) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(995) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(995);
STATE_UPDATE_MASK(996) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(996) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(996);
STATE_UPDATE_MASK(997) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(997) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(997);
STATE_UPDATE_MASK(998) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(998) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(998);
STATE_UPDATE_MASK(999) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(999) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(999);
STATE_UPDATE_MASK(1000) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1000) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1000);
STATE_UPDATE_MASK(1001) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1001) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1001);
STATE_UPDATE_MASK(1002) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1002) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1002);
STATE_UPDATE_MASK(1003) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1003) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1003);
STATE_UPDATE_MASK(1004) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1004) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1004);
STATE_UPDATE_MASK(1005) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1005) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1005);
STATE_UPDATE_MASK(1006) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1006) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1006);
STATE_UPDATE_MASK(1007) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1007) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1007);
STATE_UPDATE_MASK(1008) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1008) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1008);
STATE_UPDATE_MASK(1009) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1009) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1009);
STATE_UPDATE_MASK(1010) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1010) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1010);
STATE_UPDATE_MASK(1011) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1011) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1011);
STATE_UPDATE_MASK(1012) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1012) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1012);
STATE_UPDATE_MASK(1013) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1013) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1013);
STATE_UPDATE_MASK(1014) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1014) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1014);
STATE_UPDATE_MASK(1015) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1015) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1015);
STATE_UPDATE_MASK(1016) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1016) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1016);
STATE_UPDATE_MASK(1017) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1017) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1017);
STATE_UPDATE_MASK(1018) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1018) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1018);
STATE_UPDATE_MASK(1019) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1019) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1019);
STATE_UPDATE_MASK(1020) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1020) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1020);
STATE_UPDATE_MASK(1021) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1021) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1021);
STATE_UPDATE_MASK(1022) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1022) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1022);
STATE_UPDATE_MASK(1023) <= QEP_N_10_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1023) AND QEP_N_10_W_0_S_0_IN_CTRL_MASK(1023);

QEP_N_10_W_0_S_0_OUT_DONE <= FROM_FIRST_CU_DONE;
CONTROL_UNIT_0 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
		CONTROL_UNIT_OUT_DONE => FROM_FIRST_CU_DONE );
CONTROL_UNIT_1 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0));
CONTROL_UNIT_2 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0));
CONTROL_UNIT_3 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0));
CONTROL_UNIT_4 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_4(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_4(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_4(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_4(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_4(2 DOWNTO 0));
CONTROL_UNIT_5 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_5(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_5(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_5(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_5(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_5(2 DOWNTO 0));
CONTROL_UNIT_6 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_6(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_6(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_6(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_6(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_6(2 DOWNTO 0));
CONTROL_UNIT_7 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_7(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_7(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_7(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_7(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_7(2 DOWNTO 0));
CONTROL_UNIT_8 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_8(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_8(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_8(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_8(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_8(2 DOWNTO 0));
CONTROL_UNIT_9 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_9(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_9(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_9(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_9(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_9(2 DOWNTO 0));
CONTROL_UNIT_10 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_10(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_10(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_10(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_10(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_10(2 DOWNTO 0));
CONTROL_UNIT_11 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_11(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_11(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_11(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_11(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_11(2 DOWNTO 0));
CONTROL_UNIT_12 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_12(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_12(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_12(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_12(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_12(2 DOWNTO 0));
CONTROL_UNIT_13 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_13(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_13(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_13(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_13(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_13(2 DOWNTO 0));
CONTROL_UNIT_14 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_14(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_14(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_14(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_14(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_14(2 DOWNTO 0));
CONTROL_UNIT_15 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_15(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_15(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_15(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_15(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_15(2 DOWNTO 0));
CONTROL_UNIT_16 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_16(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_16(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_16(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_16(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_16(2 DOWNTO 0));
CONTROL_UNIT_17 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_17(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_17(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_17(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_17(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_17(2 DOWNTO 0));
CONTROL_UNIT_18 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_18(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_18(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_18(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_18(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_18(2 DOWNTO 0));
CONTROL_UNIT_19 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_19(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_19(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_19(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_19(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_19(2 DOWNTO 0));
CONTROL_UNIT_20 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_20(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_20(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_20(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_20(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_20(2 DOWNTO 0));
CONTROL_UNIT_21 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_21(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_21(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_21(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_21(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_21(2 DOWNTO 0));
CONTROL_UNIT_22 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_22(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_22(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_22(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_22(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_22(2 DOWNTO 0));
CONTROL_UNIT_23 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_23(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_23(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_23(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_23(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_23(2 DOWNTO 0));
CONTROL_UNIT_24 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_24(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_24(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_24(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_24(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_24(2 DOWNTO 0));
CONTROL_UNIT_25 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_25(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_25(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_25(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_25(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_25(2 DOWNTO 0));
CONTROL_UNIT_26 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_26(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_26(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_26(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_26(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_26(2 DOWNTO 0));
CONTROL_UNIT_27 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_27(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_27(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_27(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_27(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_27(2 DOWNTO 0));
CONTROL_UNIT_28 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_28(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_28(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_28(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_28(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_28(2 DOWNTO 0));
CONTROL_UNIT_29 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_29(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_29(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_29(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_29(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_29(2 DOWNTO 0));
CONTROL_UNIT_30 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_30(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_30(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_30(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_30(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_30(2 DOWNTO 0));
CONTROL_UNIT_31 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_31(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_31(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_31(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_31(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_31(2 DOWNTO 0));
CONTROL_UNIT_32 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_32(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_32(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_32(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_32(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_32(2 DOWNTO 0));
CONTROL_UNIT_33 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_33(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_33(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_33(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_33(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_33(2 DOWNTO 0));
CONTROL_UNIT_34 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_34(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_34(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_34(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_34(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_34(2 DOWNTO 0));
CONTROL_UNIT_35 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_35(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_35(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_35(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_35(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_35(2 DOWNTO 0));
CONTROL_UNIT_36 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_36(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_36(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_36(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_36(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_36(2 DOWNTO 0));
CONTROL_UNIT_37 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_37(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_37(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_37(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_37(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_37(2 DOWNTO 0));
CONTROL_UNIT_38 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_38(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_38(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_38(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_38(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_38(2 DOWNTO 0));
CONTROL_UNIT_39 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_39(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_39(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_39(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_39(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_39(2 DOWNTO 0));
CONTROL_UNIT_40 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_40(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_40(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_40(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_40(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_40(2 DOWNTO 0));
CONTROL_UNIT_41 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_41(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_41(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_41(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_41(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_41(2 DOWNTO 0));
CONTROL_UNIT_42 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_42(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_42(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_42(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_42(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_42(2 DOWNTO 0));
CONTROL_UNIT_43 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_43(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_43(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_43(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_43(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_43(2 DOWNTO 0));
CONTROL_UNIT_44 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_44(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_44(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_44(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_44(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_44(2 DOWNTO 0));
CONTROL_UNIT_45 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_45(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_45(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_45(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_45(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_45(2 DOWNTO 0));
CONTROL_UNIT_46 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_46(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_46(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_46(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_46(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_46(2 DOWNTO 0));
CONTROL_UNIT_47 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_47(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_47(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_47(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_47(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_47(2 DOWNTO 0));
CONTROL_UNIT_48 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_48(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_48(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_48(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_48(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_48(2 DOWNTO 0));
CONTROL_UNIT_49 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_49(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_49(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_49(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_49(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_49(2 DOWNTO 0));
CONTROL_UNIT_50 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_50(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_50(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_50(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_50(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_50(2 DOWNTO 0));
CONTROL_UNIT_51 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_51(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_51(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_51(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_51(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_51(2 DOWNTO 0));
CONTROL_UNIT_52 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_52(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_52(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_52(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_52(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_52(2 DOWNTO 0));
CONTROL_UNIT_53 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_53(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_53(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_53(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_53(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_53(2 DOWNTO 0));
CONTROL_UNIT_54 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_54(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_54(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_54(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_54(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_54(2 DOWNTO 0));
CONTROL_UNIT_55 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_55(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_55(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_55(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_55(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_55(2 DOWNTO 0));
CONTROL_UNIT_56 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_56(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_56(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_56(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_56(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_56(2 DOWNTO 0));
CONTROL_UNIT_57 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_57(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_57(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_57(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_57(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_57(2 DOWNTO 0));
CONTROL_UNIT_58 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_58(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_58(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_58(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_58(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_58(2 DOWNTO 0));
CONTROL_UNIT_59 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_59(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_59(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_59(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_59(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_59(2 DOWNTO 0));
CONTROL_UNIT_60 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_60(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_60(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_60(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_60(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_60(2 DOWNTO 0));
CONTROL_UNIT_61 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_61(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_61(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_61(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_61(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_61(2 DOWNTO 0));
CONTROL_UNIT_62 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_62(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_62(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_62(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_62(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_62(2 DOWNTO 0));
CONTROL_UNIT_63 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_63(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_63(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_63(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_63(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_63(2 DOWNTO 0));
CONTROL_UNIT_64 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_64(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_64(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_64(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_64(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_64(2 DOWNTO 0));
CONTROL_UNIT_65 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_65(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_65(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_65(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_65(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_65(2 DOWNTO 0));
CONTROL_UNIT_66 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_66(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_66(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_66(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_66(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_66(2 DOWNTO 0));
CONTROL_UNIT_67 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_67(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_67(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_67(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_67(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_67(2 DOWNTO 0));
CONTROL_UNIT_68 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_68(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_68(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_68(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_68(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_68(2 DOWNTO 0));
CONTROL_UNIT_69 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_69(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_69(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_69(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_69(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_69(2 DOWNTO 0));
CONTROL_UNIT_70 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_70(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_70(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_70(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_70(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_70(2 DOWNTO 0));
CONTROL_UNIT_71 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_71(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_71(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_71(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_71(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_71(2 DOWNTO 0));
CONTROL_UNIT_72 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_72(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_72(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_72(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_72(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_72(2 DOWNTO 0));
CONTROL_UNIT_73 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_73(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_73(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_73(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_73(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_73(2 DOWNTO 0));
CONTROL_UNIT_74 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_74(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_74(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_74(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_74(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_74(2 DOWNTO 0));
CONTROL_UNIT_75 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_75(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_75(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_75(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_75(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_75(2 DOWNTO 0));
CONTROL_UNIT_76 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_76(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_76(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_76(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_76(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_76(2 DOWNTO 0));
CONTROL_UNIT_77 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_77(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_77(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_77(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_77(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_77(2 DOWNTO 0));
CONTROL_UNIT_78 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_78(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_78(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_78(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_78(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_78(2 DOWNTO 0));
CONTROL_UNIT_79 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_79(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_79(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_79(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_79(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_79(2 DOWNTO 0));
CONTROL_UNIT_80 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_80(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_80(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_80(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_80(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_80(2 DOWNTO 0));
CONTROL_UNIT_81 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_81(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_81(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_81(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_81(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_81(2 DOWNTO 0));
CONTROL_UNIT_82 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_82(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_82(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_82(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_82(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_82(2 DOWNTO 0));
CONTROL_UNIT_83 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_83(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_83(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_83(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_83(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_83(2 DOWNTO 0));
CONTROL_UNIT_84 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_84(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_84(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_84(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_84(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_84(2 DOWNTO 0));
CONTROL_UNIT_85 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_85(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_85(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_85(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_85(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_85(2 DOWNTO 0));
CONTROL_UNIT_86 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_86(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_86(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_86(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_86(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_86(2 DOWNTO 0));
CONTROL_UNIT_87 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_87(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_87(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_87(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_87(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_87(2 DOWNTO 0));
CONTROL_UNIT_88 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_88(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_88(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_88(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_88(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_88(2 DOWNTO 0));
CONTROL_UNIT_89 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_89(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_89(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_89(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_89(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_89(2 DOWNTO 0));
CONTROL_UNIT_90 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_90(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_90(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_90(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_90(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_90(2 DOWNTO 0));
CONTROL_UNIT_91 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_91(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_91(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_91(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_91(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_91(2 DOWNTO 0));
CONTROL_UNIT_92 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_92(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_92(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_92(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_92(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_92(2 DOWNTO 0));
CONTROL_UNIT_93 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_93(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_93(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_93(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_93(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_93(2 DOWNTO 0));
CONTROL_UNIT_94 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_94(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_94(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_94(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_94(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_94(2 DOWNTO 0));
CONTROL_UNIT_95 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_95(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_95(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_95(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_95(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_95(2 DOWNTO 0));
CONTROL_UNIT_96 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_96(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_96(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_96(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_96(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_96(2 DOWNTO 0));
CONTROL_UNIT_97 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_97(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_97(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_97(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_97(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_97(2 DOWNTO 0));
CONTROL_UNIT_98 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_98(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_98(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_98(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_98(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_98(2 DOWNTO 0));
CONTROL_UNIT_99 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_99(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_99(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_99(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_99(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_99(2 DOWNTO 0));
CONTROL_UNIT_100 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_100(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_100(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_100(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_100(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_100(2 DOWNTO 0));
CONTROL_UNIT_101 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_101(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_101(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_101(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_101(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_101(2 DOWNTO 0));
CONTROL_UNIT_102 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_102(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_102(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_102(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_102(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_102(2 DOWNTO 0));
CONTROL_UNIT_103 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_103(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_103(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_103(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_103(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_103(2 DOWNTO 0));
CONTROL_UNIT_104 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_104(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_104(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_104(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_104(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_104(2 DOWNTO 0));
CONTROL_UNIT_105 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_105(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_105(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_105(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_105(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_105(2 DOWNTO 0));
CONTROL_UNIT_106 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_106(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_106(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_106(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_106(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_106(2 DOWNTO 0));
CONTROL_UNIT_107 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_107(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_107(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_107(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_107(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_107(2 DOWNTO 0));
CONTROL_UNIT_108 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_108(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_108(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_108(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_108(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_108(2 DOWNTO 0));
CONTROL_UNIT_109 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_109(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_109(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_109(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_109(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_109(2 DOWNTO 0));
CONTROL_UNIT_110 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_110(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_110(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_110(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_110(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_110(2 DOWNTO 0));
CONTROL_UNIT_111 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_111(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_111(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_111(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_111(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_111(2 DOWNTO 0));
CONTROL_UNIT_112 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_112(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_112(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_112(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_112(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_112(2 DOWNTO 0));
CONTROL_UNIT_113 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_113(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_113(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_113(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_113(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_113(2 DOWNTO 0));
CONTROL_UNIT_114 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_114(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_114(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_114(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_114(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_114(2 DOWNTO 0));
CONTROL_UNIT_115 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_115(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_115(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_115(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_115(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_115(2 DOWNTO 0));
CONTROL_UNIT_116 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_116(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_116(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_116(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_116(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_116(2 DOWNTO 0));
CONTROL_UNIT_117 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_117(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_117(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_117(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_117(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_117(2 DOWNTO 0));
CONTROL_UNIT_118 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_118(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_118(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_118(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_118(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_118(2 DOWNTO 0));
CONTROL_UNIT_119 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_119(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_119(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_119(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_119(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_119(2 DOWNTO 0));
CONTROL_UNIT_120 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_120(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_120(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_120(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_120(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_120(2 DOWNTO 0));
CONTROL_UNIT_121 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_121(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_121(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_121(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_121(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_121(2 DOWNTO 0));
CONTROL_UNIT_122 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_122(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_122(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_122(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_122(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_122(2 DOWNTO 0));
CONTROL_UNIT_123 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_123(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_123(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_123(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_123(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_123(2 DOWNTO 0));
CONTROL_UNIT_124 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_124(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_124(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_124(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_124(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_124(2 DOWNTO 0));
CONTROL_UNIT_125 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_125(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_125(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_125(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_125(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_125(2 DOWNTO 0));
CONTROL_UNIT_126 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_126(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_126(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_126(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_126(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_126(2 DOWNTO 0));
CONTROL_UNIT_127 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_127(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_127(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_127(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_127(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_127(2 DOWNTO 0));
CONTROL_UNIT_128 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_128(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_128(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_128(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_128(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_128(2 DOWNTO 0));
CONTROL_UNIT_129 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_129(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_129(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_129(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_129(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_129(2 DOWNTO 0));
CONTROL_UNIT_130 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_130(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_130(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_130(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_130(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_130(2 DOWNTO 0));
CONTROL_UNIT_131 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_131(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_131(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_131(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_131(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_131(2 DOWNTO 0));
CONTROL_UNIT_132 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_132(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_132(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_132(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_132(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_132(2 DOWNTO 0));
CONTROL_UNIT_133 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_133(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_133(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_133(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_133(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_133(2 DOWNTO 0));
CONTROL_UNIT_134 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_134(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_134(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_134(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_134(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_134(2 DOWNTO 0));
CONTROL_UNIT_135 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_135(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_135(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_135(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_135(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_135(2 DOWNTO 0));
CONTROL_UNIT_136 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_136(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_136(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_136(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_136(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_136(2 DOWNTO 0));
CONTROL_UNIT_137 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_137(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_137(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_137(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_137(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_137(2 DOWNTO 0));
CONTROL_UNIT_138 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_138(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_138(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_138(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_138(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_138(2 DOWNTO 0));
CONTROL_UNIT_139 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_139(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_139(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_139(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_139(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_139(2 DOWNTO 0));
CONTROL_UNIT_140 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_140(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_140(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_140(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_140(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_140(2 DOWNTO 0));
CONTROL_UNIT_141 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_141(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_141(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_141(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_141(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_141(2 DOWNTO 0));
CONTROL_UNIT_142 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_142(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_142(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_142(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_142(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_142(2 DOWNTO 0));
CONTROL_UNIT_143 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_143(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_143(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_143(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_143(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_143(2 DOWNTO 0));
CONTROL_UNIT_144 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_144(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_144(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_144(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_144(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_144(2 DOWNTO 0));
CONTROL_UNIT_145 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_145(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_145(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_145(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_145(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_145(2 DOWNTO 0));
CONTROL_UNIT_146 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_146(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_146(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_146(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_146(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_146(2 DOWNTO 0));
CONTROL_UNIT_147 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_147(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_147(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_147(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_147(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_147(2 DOWNTO 0));
CONTROL_UNIT_148 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_148(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_148(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_148(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_148(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_148(2 DOWNTO 0));
CONTROL_UNIT_149 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_149(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_149(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_149(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_149(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_149(2 DOWNTO 0));
CONTROL_UNIT_150 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_150(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_150(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_150(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_150(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_150(2 DOWNTO 0));
CONTROL_UNIT_151 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_151(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_151(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_151(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_151(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_151(2 DOWNTO 0));
CONTROL_UNIT_152 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_152(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_152(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_152(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_152(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_152(2 DOWNTO 0));
CONTROL_UNIT_153 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_153(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_153(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_153(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_153(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_153(2 DOWNTO 0));
CONTROL_UNIT_154 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_154(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_154(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_154(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_154(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_154(2 DOWNTO 0));
CONTROL_UNIT_155 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_155(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_155(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_155(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_155(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_155(2 DOWNTO 0));
CONTROL_UNIT_156 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_156(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_156(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_156(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_156(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_156(2 DOWNTO 0));
CONTROL_UNIT_157 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_157(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_157(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_157(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_157(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_157(2 DOWNTO 0));
CONTROL_UNIT_158 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_158(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_158(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_158(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_158(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_158(2 DOWNTO 0));
CONTROL_UNIT_159 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_159(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_159(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_159(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_159(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_159(2 DOWNTO 0));
CONTROL_UNIT_160 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_160(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_160(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_160(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_160(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_160(2 DOWNTO 0));
CONTROL_UNIT_161 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_161(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_161(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_161(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_161(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_161(2 DOWNTO 0));
CONTROL_UNIT_162 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_162(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_162(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_162(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_162(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_162(2 DOWNTO 0));
CONTROL_UNIT_163 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_163(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_163(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_163(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_163(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_163(2 DOWNTO 0));
CONTROL_UNIT_164 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_164(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_164(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_164(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_164(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_164(2 DOWNTO 0));
CONTROL_UNIT_165 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_165(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_165(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_165(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_165(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_165(2 DOWNTO 0));
CONTROL_UNIT_166 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_166(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_166(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_166(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_166(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_166(2 DOWNTO 0));
CONTROL_UNIT_167 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_167(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_167(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_167(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_167(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_167(2 DOWNTO 0));
CONTROL_UNIT_168 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_168(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_168(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_168(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_168(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_168(2 DOWNTO 0));
CONTROL_UNIT_169 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_169(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_169(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_169(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_169(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_169(2 DOWNTO 0));
CONTROL_UNIT_170 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_170(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_170(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_170(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_170(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_170(2 DOWNTO 0));
CONTROL_UNIT_171 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_171(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_171(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_171(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_171(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_171(2 DOWNTO 0));
CONTROL_UNIT_172 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_172(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_172(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_172(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_172(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_172(2 DOWNTO 0));
CONTROL_UNIT_173 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_173(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_173(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_173(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_173(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_173(2 DOWNTO 0));
CONTROL_UNIT_174 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_174(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_174(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_174(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_174(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_174(2 DOWNTO 0));
CONTROL_UNIT_175 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_175(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_175(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_175(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_175(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_175(2 DOWNTO 0));
CONTROL_UNIT_176 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_176(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_176(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_176(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_176(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_176(2 DOWNTO 0));
CONTROL_UNIT_177 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_177(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_177(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_177(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_177(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_177(2 DOWNTO 0));
CONTROL_UNIT_178 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_178(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_178(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_178(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_178(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_178(2 DOWNTO 0));
CONTROL_UNIT_179 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_179(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_179(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_179(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_179(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_179(2 DOWNTO 0));
CONTROL_UNIT_180 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_180(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_180(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_180(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_180(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_180(2 DOWNTO 0));
CONTROL_UNIT_181 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_181(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_181(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_181(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_181(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_181(2 DOWNTO 0));
CONTROL_UNIT_182 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_182(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_182(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_182(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_182(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_182(2 DOWNTO 0));
CONTROL_UNIT_183 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_183(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_183(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_183(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_183(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_183(2 DOWNTO 0));
CONTROL_UNIT_184 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_184(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_184(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_184(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_184(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_184(2 DOWNTO 0));
CONTROL_UNIT_185 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_185(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_185(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_185(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_185(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_185(2 DOWNTO 0));
CONTROL_UNIT_186 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_186(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_186(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_186(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_186(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_186(2 DOWNTO 0));
CONTROL_UNIT_187 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_187(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_187(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_187(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_187(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_187(2 DOWNTO 0));
CONTROL_UNIT_188 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_188(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_188(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_188(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_188(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_188(2 DOWNTO 0));
CONTROL_UNIT_189 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_189(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_189(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_189(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_189(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_189(2 DOWNTO 0));
CONTROL_UNIT_190 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_190(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_190(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_190(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_190(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_190(2 DOWNTO 0));
CONTROL_UNIT_191 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_191(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_191(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_191(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_191(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_191(2 DOWNTO 0));
CONTROL_UNIT_192 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_192(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_192(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_192(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_192(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_192(2 DOWNTO 0));
CONTROL_UNIT_193 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_193(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_193(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_193(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_193(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_193(2 DOWNTO 0));
CONTROL_UNIT_194 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_194(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_194(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_194(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_194(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_194(2 DOWNTO 0));
CONTROL_UNIT_195 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_195(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_195(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_195(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_195(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_195(2 DOWNTO 0));
CONTROL_UNIT_196 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_196(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_196(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_196(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_196(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_196(2 DOWNTO 0));
CONTROL_UNIT_197 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_197(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_197(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_197(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_197(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_197(2 DOWNTO 0));
CONTROL_UNIT_198 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_198(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_198(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_198(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_198(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_198(2 DOWNTO 0));
CONTROL_UNIT_199 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_199(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_199(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_199(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_199(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_199(2 DOWNTO 0));
CONTROL_UNIT_200 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_200(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_200(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_200(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_200(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_200(2 DOWNTO 0));
CONTROL_UNIT_201 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_201(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_201(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_201(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_201(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_201(2 DOWNTO 0));
CONTROL_UNIT_202 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_202(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_202(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_202(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_202(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_202(2 DOWNTO 0));
CONTROL_UNIT_203 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_203(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_203(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_203(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_203(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_203(2 DOWNTO 0));
CONTROL_UNIT_204 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_204(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_204(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_204(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_204(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_204(2 DOWNTO 0));
CONTROL_UNIT_205 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_205(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_205(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_205(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_205(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_205(2 DOWNTO 0));
CONTROL_UNIT_206 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_206(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_206(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_206(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_206(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_206(2 DOWNTO 0));
CONTROL_UNIT_207 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_207(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_207(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_207(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_207(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_207(2 DOWNTO 0));
CONTROL_UNIT_208 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_208(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_208(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_208(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_208(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_208(2 DOWNTO 0));
CONTROL_UNIT_209 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_209(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_209(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_209(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_209(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_209(2 DOWNTO 0));
CONTROL_UNIT_210 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_210(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_210(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_210(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_210(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_210(2 DOWNTO 0));
CONTROL_UNIT_211 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_211(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_211(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_211(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_211(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_211(2 DOWNTO 0));
CONTROL_UNIT_212 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_212(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_212(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_212(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_212(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_212(2 DOWNTO 0));
CONTROL_UNIT_213 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_213(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_213(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_213(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_213(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_213(2 DOWNTO 0));
CONTROL_UNIT_214 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_214(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_214(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_214(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_214(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_214(2 DOWNTO 0));
CONTROL_UNIT_215 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_215(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_215(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_215(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_215(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_215(2 DOWNTO 0));
CONTROL_UNIT_216 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_216(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_216(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_216(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_216(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_216(2 DOWNTO 0));
CONTROL_UNIT_217 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_217(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_217(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_217(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_217(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_217(2 DOWNTO 0));
CONTROL_UNIT_218 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_218(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_218(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_218(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_218(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_218(2 DOWNTO 0));
CONTROL_UNIT_219 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_219(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_219(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_219(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_219(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_219(2 DOWNTO 0));
CONTROL_UNIT_220 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_220(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_220(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_220(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_220(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_220(2 DOWNTO 0));
CONTROL_UNIT_221 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_221(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_221(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_221(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_221(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_221(2 DOWNTO 0));
CONTROL_UNIT_222 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_222(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_222(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_222(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_222(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_222(2 DOWNTO 0));
CONTROL_UNIT_223 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_223(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_223(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_223(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_223(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_223(2 DOWNTO 0));
CONTROL_UNIT_224 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_224(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_224(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_224(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_224(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_224(2 DOWNTO 0));
CONTROL_UNIT_225 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_225(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_225(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_225(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_225(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_225(2 DOWNTO 0));
CONTROL_UNIT_226 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_226(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_226(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_226(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_226(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_226(2 DOWNTO 0));
CONTROL_UNIT_227 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_227(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_227(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_227(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_227(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_227(2 DOWNTO 0));
CONTROL_UNIT_228 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_228(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_228(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_228(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_228(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_228(2 DOWNTO 0));
CONTROL_UNIT_229 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_229(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_229(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_229(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_229(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_229(2 DOWNTO 0));
CONTROL_UNIT_230 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_230(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_230(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_230(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_230(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_230(2 DOWNTO 0));
CONTROL_UNIT_231 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_231(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_231(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_231(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_231(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_231(2 DOWNTO 0));
CONTROL_UNIT_232 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_232(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_232(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_232(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_232(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_232(2 DOWNTO 0));
CONTROL_UNIT_233 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_233(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_233(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_233(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_233(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_233(2 DOWNTO 0));
CONTROL_UNIT_234 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_234(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_234(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_234(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_234(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_234(2 DOWNTO 0));
CONTROL_UNIT_235 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_235(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_235(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_235(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_235(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_235(2 DOWNTO 0));
CONTROL_UNIT_236 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_236(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_236(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_236(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_236(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_236(2 DOWNTO 0));
CONTROL_UNIT_237 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_237(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_237(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_237(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_237(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_237(2 DOWNTO 0));
CONTROL_UNIT_238 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_238(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_238(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_238(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_238(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_238(2 DOWNTO 0));
CONTROL_UNIT_239 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_239(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_239(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_239(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_239(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_239(2 DOWNTO 0));
CONTROL_UNIT_240 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_240(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_240(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_240(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_240(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_240(2 DOWNTO 0));
CONTROL_UNIT_241 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_241(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_241(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_241(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_241(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_241(2 DOWNTO 0));
CONTROL_UNIT_242 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_242(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_242(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_242(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_242(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_242(2 DOWNTO 0));
CONTROL_UNIT_243 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_243(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_243(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_243(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_243(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_243(2 DOWNTO 0));
CONTROL_UNIT_244 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_244(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_244(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_244(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_244(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_244(2 DOWNTO 0));
CONTROL_UNIT_245 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_245(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_245(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_245(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_245(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_245(2 DOWNTO 0));
CONTROL_UNIT_246 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_246(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_246(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_246(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_246(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_246(2 DOWNTO 0));
CONTROL_UNIT_247 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_247(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_247(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_247(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_247(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_247(2 DOWNTO 0));
CONTROL_UNIT_248 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_248(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_248(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_248(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_248(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_248(2 DOWNTO 0));
CONTROL_UNIT_249 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_249(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_249(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_249(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_249(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_249(2 DOWNTO 0));
CONTROL_UNIT_250 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_250(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_250(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_250(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_250(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_250(2 DOWNTO 0));
CONTROL_UNIT_251 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_251(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_251(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_251(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_251(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_251(2 DOWNTO 0));
CONTROL_UNIT_252 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_252(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_252(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_252(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_252(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_252(2 DOWNTO 0));
CONTROL_UNIT_253 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_253(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_253(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_253(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_253(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_253(2 DOWNTO 0));
CONTROL_UNIT_254 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_254(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_254(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_254(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_254(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_254(2 DOWNTO 0));
CONTROL_UNIT_255 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_255(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_255(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_255(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_255(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_255(2 DOWNTO 0));
CONTROL_UNIT_256 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_256(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_256(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_256(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_256(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_256(2 DOWNTO 0));
CONTROL_UNIT_257 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_257(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_257(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_257(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_257(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_257(2 DOWNTO 0));
CONTROL_UNIT_258 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_258(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_258(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_258(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_258(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_258(2 DOWNTO 0));
CONTROL_UNIT_259 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_259(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_259(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_259(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_259(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_259(2 DOWNTO 0));
CONTROL_UNIT_260 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_260(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_260(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_260(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_260(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_260(2 DOWNTO 0));
CONTROL_UNIT_261 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_261(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_261(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_261(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_261(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_261(2 DOWNTO 0));
CONTROL_UNIT_262 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_262(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_262(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_262(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_262(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_262(2 DOWNTO 0));
CONTROL_UNIT_263 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_263(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_263(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_263(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_263(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_263(2 DOWNTO 0));
CONTROL_UNIT_264 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_264(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_264(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_264(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_264(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_264(2 DOWNTO 0));
CONTROL_UNIT_265 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_265(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_265(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_265(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_265(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_265(2 DOWNTO 0));
CONTROL_UNIT_266 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_266(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_266(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_266(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_266(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_266(2 DOWNTO 0));
CONTROL_UNIT_267 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_267(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_267(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_267(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_267(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_267(2 DOWNTO 0));
CONTROL_UNIT_268 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_268(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_268(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_268(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_268(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_268(2 DOWNTO 0));
CONTROL_UNIT_269 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_269(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_269(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_269(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_269(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_269(2 DOWNTO 0));
CONTROL_UNIT_270 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_270(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_270(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_270(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_270(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_270(2 DOWNTO 0));
CONTROL_UNIT_271 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_271(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_271(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_271(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_271(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_271(2 DOWNTO 0));
CONTROL_UNIT_272 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_272(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_272(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_272(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_272(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_272(2 DOWNTO 0));
CONTROL_UNIT_273 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_273(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_273(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_273(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_273(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_273(2 DOWNTO 0));
CONTROL_UNIT_274 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_274(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_274(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_274(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_274(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_274(2 DOWNTO 0));
CONTROL_UNIT_275 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_275(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_275(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_275(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_275(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_275(2 DOWNTO 0));
CONTROL_UNIT_276 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_276(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_276(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_276(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_276(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_276(2 DOWNTO 0));
CONTROL_UNIT_277 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_277(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_277(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_277(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_277(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_277(2 DOWNTO 0));
CONTROL_UNIT_278 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_278(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_278(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_278(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_278(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_278(2 DOWNTO 0));
CONTROL_UNIT_279 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_279(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_279(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_279(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_279(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_279(2 DOWNTO 0));
CONTROL_UNIT_280 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_280(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_280(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_280(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_280(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_280(2 DOWNTO 0));
CONTROL_UNIT_281 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_281(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_281(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_281(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_281(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_281(2 DOWNTO 0));
CONTROL_UNIT_282 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_282(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_282(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_282(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_282(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_282(2 DOWNTO 0));
CONTROL_UNIT_283 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_283(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_283(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_283(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_283(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_283(2 DOWNTO 0));
CONTROL_UNIT_284 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_284(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_284(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_284(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_284(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_284(2 DOWNTO 0));
CONTROL_UNIT_285 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_285(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_285(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_285(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_285(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_285(2 DOWNTO 0));
CONTROL_UNIT_286 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_286(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_286(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_286(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_286(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_286(2 DOWNTO 0));
CONTROL_UNIT_287 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_287(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_287(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_287(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_287(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_287(2 DOWNTO 0));
CONTROL_UNIT_288 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_288(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_288(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_288(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_288(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_288(2 DOWNTO 0));
CONTROL_UNIT_289 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_289(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_289(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_289(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_289(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_289(2 DOWNTO 0));
CONTROL_UNIT_290 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_290(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_290(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_290(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_290(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_290(2 DOWNTO 0));
CONTROL_UNIT_291 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_291(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_291(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_291(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_291(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_291(2 DOWNTO 0));
CONTROL_UNIT_292 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_292(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_292(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_292(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_292(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_292(2 DOWNTO 0));
CONTROL_UNIT_293 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_293(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_293(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_293(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_293(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_293(2 DOWNTO 0));
CONTROL_UNIT_294 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_294(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_294(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_294(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_294(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_294(2 DOWNTO 0));
CONTROL_UNIT_295 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_295(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_295(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_295(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_295(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_295(2 DOWNTO 0));
CONTROL_UNIT_296 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_296(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_296(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_296(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_296(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_296(2 DOWNTO 0));
CONTROL_UNIT_297 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_297(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_297(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_297(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_297(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_297(2 DOWNTO 0));
CONTROL_UNIT_298 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_298(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_298(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_298(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_298(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_298(2 DOWNTO 0));
CONTROL_UNIT_299 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_299(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_299(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_299(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_299(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_299(2 DOWNTO 0));
CONTROL_UNIT_300 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_300(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_300(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_300(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_300(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_300(2 DOWNTO 0));
CONTROL_UNIT_301 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_301(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_301(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_301(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_301(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_301(2 DOWNTO 0));
CONTROL_UNIT_302 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_302(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_302(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_302(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_302(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_302(2 DOWNTO 0));
CONTROL_UNIT_303 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_303(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_303(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_303(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_303(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_303(2 DOWNTO 0));
CONTROL_UNIT_304 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_304(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_304(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_304(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_304(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_304(2 DOWNTO 0));
CONTROL_UNIT_305 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_305(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_305(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_305(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_305(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_305(2 DOWNTO 0));
CONTROL_UNIT_306 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_306(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_306(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_306(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_306(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_306(2 DOWNTO 0));
CONTROL_UNIT_307 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_307(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_307(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_307(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_307(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_307(2 DOWNTO 0));
CONTROL_UNIT_308 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_308(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_308(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_308(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_308(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_308(2 DOWNTO 0));
CONTROL_UNIT_309 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_309(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_309(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_309(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_309(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_309(2 DOWNTO 0));
CONTROL_UNIT_310 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_310(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_310(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_310(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_310(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_310(2 DOWNTO 0));
CONTROL_UNIT_311 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_311(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_311(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_311(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_311(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_311(2 DOWNTO 0));
CONTROL_UNIT_312 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_312(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_312(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_312(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_312(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_312(2 DOWNTO 0));
CONTROL_UNIT_313 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_313(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_313(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_313(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_313(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_313(2 DOWNTO 0));
CONTROL_UNIT_314 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_314(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_314(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_314(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_314(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_314(2 DOWNTO 0));
CONTROL_UNIT_315 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_315(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_315(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_315(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_315(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_315(2 DOWNTO 0));
CONTROL_UNIT_316 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_316(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_316(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_316(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_316(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_316(2 DOWNTO 0));
CONTROL_UNIT_317 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_317(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_317(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_317(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_317(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_317(2 DOWNTO 0));
CONTROL_UNIT_318 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_318(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_318(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_318(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_318(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_318(2 DOWNTO 0));
CONTROL_UNIT_319 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_319(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_319(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_319(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_319(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_319(2 DOWNTO 0));
CONTROL_UNIT_320 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_320(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_320(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_320(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_320(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_320(2 DOWNTO 0));
CONTROL_UNIT_321 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_321(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_321(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_321(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_321(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_321(2 DOWNTO 0));
CONTROL_UNIT_322 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_322(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_322(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_322(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_322(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_322(2 DOWNTO 0));
CONTROL_UNIT_323 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_323(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_323(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_323(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_323(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_323(2 DOWNTO 0));
CONTROL_UNIT_324 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_324(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_324(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_324(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_324(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_324(2 DOWNTO 0));
CONTROL_UNIT_325 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_325(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_325(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_325(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_325(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_325(2 DOWNTO 0));
CONTROL_UNIT_326 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_326(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_326(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_326(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_326(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_326(2 DOWNTO 0));
CONTROL_UNIT_327 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_327(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_327(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_327(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_327(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_327(2 DOWNTO 0));
CONTROL_UNIT_328 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_328(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_328(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_328(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_328(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_328(2 DOWNTO 0));
CONTROL_UNIT_329 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_329(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_329(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_329(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_329(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_329(2 DOWNTO 0));
CONTROL_UNIT_330 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_330(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_330(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_330(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_330(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_330(2 DOWNTO 0));
CONTROL_UNIT_331 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_331(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_331(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_331(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_331(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_331(2 DOWNTO 0));
CONTROL_UNIT_332 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_332(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_332(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_332(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_332(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_332(2 DOWNTO 0));
CONTROL_UNIT_333 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_333(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_333(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_333(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_333(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_333(2 DOWNTO 0));
CONTROL_UNIT_334 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_334(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_334(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_334(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_334(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_334(2 DOWNTO 0));
CONTROL_UNIT_335 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_335(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_335(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_335(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_335(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_335(2 DOWNTO 0));
CONTROL_UNIT_336 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_336(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_336(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_336(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_336(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_336(2 DOWNTO 0));
CONTROL_UNIT_337 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_337(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_337(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_337(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_337(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_337(2 DOWNTO 0));
CONTROL_UNIT_338 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_338(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_338(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_338(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_338(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_338(2 DOWNTO 0));
CONTROL_UNIT_339 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_339(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_339(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_339(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_339(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_339(2 DOWNTO 0));
CONTROL_UNIT_340 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_340(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_340(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_340(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_340(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_340(2 DOWNTO 0));
CONTROL_UNIT_341 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_341(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_341(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_341(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_341(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_341(2 DOWNTO 0));
CONTROL_UNIT_342 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_342(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_342(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_342(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_342(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_342(2 DOWNTO 0));
CONTROL_UNIT_343 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_343(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_343(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_343(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_343(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_343(2 DOWNTO 0));
CONTROL_UNIT_344 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_344(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_344(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_344(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_344(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_344(2 DOWNTO 0));
CONTROL_UNIT_345 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_345(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_345(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_345(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_345(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_345(2 DOWNTO 0));
CONTROL_UNIT_346 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_346(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_346(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_346(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_346(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_346(2 DOWNTO 0));
CONTROL_UNIT_347 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_347(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_347(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_347(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_347(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_347(2 DOWNTO 0));
CONTROL_UNIT_348 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_348(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_348(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_348(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_348(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_348(2 DOWNTO 0));
CONTROL_UNIT_349 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_349(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_349(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_349(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_349(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_349(2 DOWNTO 0));
CONTROL_UNIT_350 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_350(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_350(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_350(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_350(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_350(2 DOWNTO 0));
CONTROL_UNIT_351 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_351(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_351(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_351(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_351(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_351(2 DOWNTO 0));
CONTROL_UNIT_352 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_352(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_352(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_352(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_352(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_352(2 DOWNTO 0));
CONTROL_UNIT_353 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_353(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_353(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_353(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_353(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_353(2 DOWNTO 0));
CONTROL_UNIT_354 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_354(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_354(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_354(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_354(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_354(2 DOWNTO 0));
CONTROL_UNIT_355 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_355(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_355(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_355(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_355(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_355(2 DOWNTO 0));
CONTROL_UNIT_356 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_356(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_356(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_356(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_356(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_356(2 DOWNTO 0));
CONTROL_UNIT_357 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_357(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_357(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_357(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_357(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_357(2 DOWNTO 0));
CONTROL_UNIT_358 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_358(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_358(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_358(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_358(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_358(2 DOWNTO 0));
CONTROL_UNIT_359 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_359(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_359(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_359(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_359(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_359(2 DOWNTO 0));
CONTROL_UNIT_360 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_360(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_360(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_360(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_360(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_360(2 DOWNTO 0));
CONTROL_UNIT_361 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_361(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_361(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_361(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_361(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_361(2 DOWNTO 0));
CONTROL_UNIT_362 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_362(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_362(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_362(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_362(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_362(2 DOWNTO 0));
CONTROL_UNIT_363 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_363(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_363(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_363(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_363(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_363(2 DOWNTO 0));
CONTROL_UNIT_364 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_364(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_364(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_364(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_364(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_364(2 DOWNTO 0));
CONTROL_UNIT_365 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_365(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_365(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_365(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_365(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_365(2 DOWNTO 0));
CONTROL_UNIT_366 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_366(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_366(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_366(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_366(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_366(2 DOWNTO 0));
CONTROL_UNIT_367 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_367(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_367(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_367(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_367(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_367(2 DOWNTO 0));
CONTROL_UNIT_368 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_368(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_368(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_368(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_368(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_368(2 DOWNTO 0));
CONTROL_UNIT_369 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_369(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_369(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_369(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_369(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_369(2 DOWNTO 0));
CONTROL_UNIT_370 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_370(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_370(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_370(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_370(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_370(2 DOWNTO 0));
CONTROL_UNIT_371 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_371(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_371(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_371(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_371(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_371(2 DOWNTO 0));
CONTROL_UNIT_372 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_372(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_372(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_372(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_372(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_372(2 DOWNTO 0));
CONTROL_UNIT_373 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_373(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_373(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_373(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_373(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_373(2 DOWNTO 0));
CONTROL_UNIT_374 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_374(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_374(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_374(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_374(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_374(2 DOWNTO 0));
CONTROL_UNIT_375 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_375(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_375(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_375(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_375(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_375(2 DOWNTO 0));
CONTROL_UNIT_376 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_376(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_376(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_376(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_376(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_376(2 DOWNTO 0));
CONTROL_UNIT_377 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_377(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_377(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_377(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_377(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_377(2 DOWNTO 0));
CONTROL_UNIT_378 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_378(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_378(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_378(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_378(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_378(2 DOWNTO 0));
CONTROL_UNIT_379 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_379(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_379(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_379(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_379(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_379(2 DOWNTO 0));
CONTROL_UNIT_380 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_380(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_380(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_380(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_380(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_380(2 DOWNTO 0));
CONTROL_UNIT_381 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_381(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_381(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_381(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_381(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_381(2 DOWNTO 0));
CONTROL_UNIT_382 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_382(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_382(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_382(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_382(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_382(2 DOWNTO 0));
CONTROL_UNIT_383 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_383(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_383(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_383(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_383(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_383(2 DOWNTO 0));
CONTROL_UNIT_384 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_384(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_384(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_384(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_384(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_384(2 DOWNTO 0));
CONTROL_UNIT_385 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_385(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_385(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_385(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_385(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_385(2 DOWNTO 0));
CONTROL_UNIT_386 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_386(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_386(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_386(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_386(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_386(2 DOWNTO 0));
CONTROL_UNIT_387 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_387(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_387(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_387(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_387(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_387(2 DOWNTO 0));
CONTROL_UNIT_388 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_388(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_388(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_388(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_388(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_388(2 DOWNTO 0));
CONTROL_UNIT_389 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_389(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_389(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_389(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_389(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_389(2 DOWNTO 0));
CONTROL_UNIT_390 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_390(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_390(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_390(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_390(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_390(2 DOWNTO 0));
CONTROL_UNIT_391 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_391(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_391(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_391(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_391(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_391(2 DOWNTO 0));
CONTROL_UNIT_392 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_392(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_392(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_392(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_392(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_392(2 DOWNTO 0));
CONTROL_UNIT_393 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_393(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_393(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_393(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_393(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_393(2 DOWNTO 0));
CONTROL_UNIT_394 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_394(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_394(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_394(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_394(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_394(2 DOWNTO 0));
CONTROL_UNIT_395 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_395(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_395(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_395(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_395(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_395(2 DOWNTO 0));
CONTROL_UNIT_396 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_396(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_396(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_396(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_396(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_396(2 DOWNTO 0));
CONTROL_UNIT_397 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_397(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_397(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_397(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_397(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_397(2 DOWNTO 0));
CONTROL_UNIT_398 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_398(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_398(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_398(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_398(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_398(2 DOWNTO 0));
CONTROL_UNIT_399 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_399(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_399(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_399(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_399(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_399(2 DOWNTO 0));
CONTROL_UNIT_400 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_400(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_400(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_400(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_400(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_400(2 DOWNTO 0));
CONTROL_UNIT_401 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_401(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_401(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_401(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_401(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_401(2 DOWNTO 0));
CONTROL_UNIT_402 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_402(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_402(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_402(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_402(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_402(2 DOWNTO 0));
CONTROL_UNIT_403 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_403(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_403(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_403(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_403(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_403(2 DOWNTO 0));
CONTROL_UNIT_404 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_404(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_404(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_404(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_404(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_404(2 DOWNTO 0));
CONTROL_UNIT_405 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_405(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_405(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_405(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_405(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_405(2 DOWNTO 0));
CONTROL_UNIT_406 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_406(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_406(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_406(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_406(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_406(2 DOWNTO 0));
CONTROL_UNIT_407 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_407(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_407(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_407(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_407(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_407(2 DOWNTO 0));
CONTROL_UNIT_408 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_408(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_408(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_408(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_408(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_408(2 DOWNTO 0));
CONTROL_UNIT_409 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_409(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_409(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_409(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_409(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_409(2 DOWNTO 0));
CONTROL_UNIT_410 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_410(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_410(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_410(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_410(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_410(2 DOWNTO 0));
CONTROL_UNIT_411 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_411(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_411(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_411(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_411(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_411(2 DOWNTO 0));
CONTROL_UNIT_412 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_412(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_412(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_412(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_412(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_412(2 DOWNTO 0));
CONTROL_UNIT_413 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_413(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_413(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_413(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_413(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_413(2 DOWNTO 0));
CONTROL_UNIT_414 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_414(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_414(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_414(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_414(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_414(2 DOWNTO 0));
CONTROL_UNIT_415 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_415(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_415(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_415(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_415(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_415(2 DOWNTO 0));
CONTROL_UNIT_416 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_416(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_416(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_416(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_416(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_416(2 DOWNTO 0));
CONTROL_UNIT_417 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_417(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_417(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_417(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_417(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_417(2 DOWNTO 0));
CONTROL_UNIT_418 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_418(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_418(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_418(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_418(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_418(2 DOWNTO 0));
CONTROL_UNIT_419 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_419(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_419(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_419(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_419(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_419(2 DOWNTO 0));
CONTROL_UNIT_420 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_420(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_420(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_420(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_420(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_420(2 DOWNTO 0));
CONTROL_UNIT_421 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_421(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_421(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_421(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_421(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_421(2 DOWNTO 0));
CONTROL_UNIT_422 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_422(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_422(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_422(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_422(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_422(2 DOWNTO 0));
CONTROL_UNIT_423 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_423(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_423(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_423(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_423(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_423(2 DOWNTO 0));
CONTROL_UNIT_424 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_424(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_424(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_424(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_424(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_424(2 DOWNTO 0));
CONTROL_UNIT_425 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_425(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_425(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_425(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_425(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_425(2 DOWNTO 0));
CONTROL_UNIT_426 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_426(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_426(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_426(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_426(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_426(2 DOWNTO 0));
CONTROL_UNIT_427 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_427(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_427(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_427(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_427(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_427(2 DOWNTO 0));
CONTROL_UNIT_428 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_428(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_428(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_428(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_428(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_428(2 DOWNTO 0));
CONTROL_UNIT_429 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_429(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_429(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_429(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_429(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_429(2 DOWNTO 0));
CONTROL_UNIT_430 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_430(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_430(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_430(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_430(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_430(2 DOWNTO 0));
CONTROL_UNIT_431 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_431(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_431(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_431(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_431(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_431(2 DOWNTO 0));
CONTROL_UNIT_432 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_432(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_432(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_432(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_432(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_432(2 DOWNTO 0));
CONTROL_UNIT_433 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_433(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_433(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_433(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_433(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_433(2 DOWNTO 0));
CONTROL_UNIT_434 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_434(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_434(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_434(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_434(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_434(2 DOWNTO 0));
CONTROL_UNIT_435 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_435(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_435(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_435(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_435(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_435(2 DOWNTO 0));
CONTROL_UNIT_436 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_436(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_436(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_436(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_436(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_436(2 DOWNTO 0));
CONTROL_UNIT_437 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_437(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_437(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_437(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_437(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_437(2 DOWNTO 0));
CONTROL_UNIT_438 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_438(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_438(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_438(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_438(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_438(2 DOWNTO 0));
CONTROL_UNIT_439 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_439(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_439(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_439(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_439(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_439(2 DOWNTO 0));
CONTROL_UNIT_440 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_440(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_440(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_440(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_440(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_440(2 DOWNTO 0));
CONTROL_UNIT_441 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_441(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_441(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_441(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_441(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_441(2 DOWNTO 0));
CONTROL_UNIT_442 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_442(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_442(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_442(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_442(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_442(2 DOWNTO 0));
CONTROL_UNIT_443 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_443(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_443(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_443(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_443(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_443(2 DOWNTO 0));
CONTROL_UNIT_444 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_444(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_444(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_444(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_444(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_444(2 DOWNTO 0));
CONTROL_UNIT_445 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_445(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_445(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_445(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_445(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_445(2 DOWNTO 0));
CONTROL_UNIT_446 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_446(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_446(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_446(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_446(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_446(2 DOWNTO 0));
CONTROL_UNIT_447 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_447(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_447(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_447(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_447(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_447(2 DOWNTO 0));
CONTROL_UNIT_448 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_448(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_448(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_448(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_448(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_448(2 DOWNTO 0));
CONTROL_UNIT_449 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_449(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_449(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_449(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_449(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_449(2 DOWNTO 0));
CONTROL_UNIT_450 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_450(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_450(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_450(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_450(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_450(2 DOWNTO 0));
CONTROL_UNIT_451 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_451(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_451(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_451(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_451(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_451(2 DOWNTO 0));
CONTROL_UNIT_452 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_452(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_452(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_452(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_452(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_452(2 DOWNTO 0));
CONTROL_UNIT_453 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_453(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_453(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_453(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_453(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_453(2 DOWNTO 0));
CONTROL_UNIT_454 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_454(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_454(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_454(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_454(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_454(2 DOWNTO 0));
CONTROL_UNIT_455 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_455(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_455(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_455(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_455(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_455(2 DOWNTO 0));
CONTROL_UNIT_456 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_456(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_456(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_456(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_456(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_456(2 DOWNTO 0));
CONTROL_UNIT_457 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_457(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_457(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_457(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_457(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_457(2 DOWNTO 0));
CONTROL_UNIT_458 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_458(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_458(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_458(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_458(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_458(2 DOWNTO 0));
CONTROL_UNIT_459 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_459(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_459(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_459(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_459(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_459(2 DOWNTO 0));
CONTROL_UNIT_460 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_460(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_460(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_460(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_460(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_460(2 DOWNTO 0));
CONTROL_UNIT_461 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_461(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_461(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_461(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_461(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_461(2 DOWNTO 0));
CONTROL_UNIT_462 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_462(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_462(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_462(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_462(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_462(2 DOWNTO 0));
CONTROL_UNIT_463 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_463(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_463(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_463(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_463(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_463(2 DOWNTO 0));
CONTROL_UNIT_464 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_464(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_464(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_464(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_464(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_464(2 DOWNTO 0));
CONTROL_UNIT_465 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_465(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_465(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_465(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_465(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_465(2 DOWNTO 0));
CONTROL_UNIT_466 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_466(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_466(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_466(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_466(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_466(2 DOWNTO 0));
CONTROL_UNIT_467 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_467(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_467(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_467(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_467(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_467(2 DOWNTO 0));
CONTROL_UNIT_468 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_468(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_468(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_468(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_468(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_468(2 DOWNTO 0));
CONTROL_UNIT_469 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_469(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_469(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_469(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_469(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_469(2 DOWNTO 0));
CONTROL_UNIT_470 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_470(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_470(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_470(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_470(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_470(2 DOWNTO 0));
CONTROL_UNIT_471 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_471(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_471(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_471(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_471(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_471(2 DOWNTO 0));
CONTROL_UNIT_472 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_472(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_472(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_472(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_472(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_472(2 DOWNTO 0));
CONTROL_UNIT_473 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_473(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_473(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_473(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_473(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_473(2 DOWNTO 0));
CONTROL_UNIT_474 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_474(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_474(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_474(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_474(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_474(2 DOWNTO 0));
CONTROL_UNIT_475 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_475(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_475(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_475(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_475(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_475(2 DOWNTO 0));
CONTROL_UNIT_476 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_476(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_476(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_476(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_476(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_476(2 DOWNTO 0));
CONTROL_UNIT_477 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_477(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_477(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_477(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_477(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_477(2 DOWNTO 0));
CONTROL_UNIT_478 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_478(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_478(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_478(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_478(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_478(2 DOWNTO 0));
CONTROL_UNIT_479 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_479(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_479(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_479(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_479(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_479(2 DOWNTO 0));
CONTROL_UNIT_480 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_480(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_480(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_480(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_480(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_480(2 DOWNTO 0));
CONTROL_UNIT_481 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_481(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_481(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_481(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_481(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_481(2 DOWNTO 0));
CONTROL_UNIT_482 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_482(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_482(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_482(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_482(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_482(2 DOWNTO 0));
CONTROL_UNIT_483 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_483(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_483(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_483(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_483(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_483(2 DOWNTO 0));
CONTROL_UNIT_484 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_484(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_484(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_484(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_484(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_484(2 DOWNTO 0));
CONTROL_UNIT_485 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_485(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_485(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_485(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_485(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_485(2 DOWNTO 0));
CONTROL_UNIT_486 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_486(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_486(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_486(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_486(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_486(2 DOWNTO 0));
CONTROL_UNIT_487 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_487(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_487(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_487(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_487(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_487(2 DOWNTO 0));
CONTROL_UNIT_488 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_488(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_488(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_488(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_488(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_488(2 DOWNTO 0));
CONTROL_UNIT_489 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_489(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_489(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_489(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_489(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_489(2 DOWNTO 0));
CONTROL_UNIT_490 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_490(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_490(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_490(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_490(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_490(2 DOWNTO 0));
CONTROL_UNIT_491 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_491(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_491(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_491(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_491(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_491(2 DOWNTO 0));
CONTROL_UNIT_492 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_492(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_492(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_492(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_492(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_492(2 DOWNTO 0));
CONTROL_UNIT_493 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_493(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_493(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_493(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_493(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_493(2 DOWNTO 0));
CONTROL_UNIT_494 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_494(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_494(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_494(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_494(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_494(2 DOWNTO 0));
CONTROL_UNIT_495 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_495(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_495(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_495(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_495(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_495(2 DOWNTO 0));
CONTROL_UNIT_496 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_496(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_496(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_496(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_496(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_496(2 DOWNTO 0));
CONTROL_UNIT_497 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_497(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_497(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_497(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_497(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_497(2 DOWNTO 0));
CONTROL_UNIT_498 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_498(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_498(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_498(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_498(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_498(2 DOWNTO 0));
CONTROL_UNIT_499 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_499(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_499(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_499(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_499(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_499(2 DOWNTO 0));
CONTROL_UNIT_500 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_500(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_500(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_500(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_500(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_500(2 DOWNTO 0));
CONTROL_UNIT_501 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_501(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_501(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_501(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_501(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_501(2 DOWNTO 0));
CONTROL_UNIT_502 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_502(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_502(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_502(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_502(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_502(2 DOWNTO 0));
CONTROL_UNIT_503 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_503(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_503(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_503(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_503(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_503(2 DOWNTO 0));
CONTROL_UNIT_504 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_504(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_504(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_504(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_504(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_504(2 DOWNTO 0));
CONTROL_UNIT_505 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_505(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_505(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_505(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_505(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_505(2 DOWNTO 0));
CONTROL_UNIT_506 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_506(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_506(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_506(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_506(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_506(2 DOWNTO 0));
CONTROL_UNIT_507 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_507(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_507(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_507(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_507(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_507(2 DOWNTO 0));
CONTROL_UNIT_508 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_508(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_508(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_508(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_508(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_508(2 DOWNTO 0));
CONTROL_UNIT_509 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_509(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_509(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_509(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_509(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_509(2 DOWNTO 0));
CONTROL_UNIT_510 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_510(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_510(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_510(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_510(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_510(2 DOWNTO 0));
CONTROL_UNIT_511 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_10_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_10_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_511(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_511(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_511(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_511(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_511(2 DOWNTO 0));

DATAPATH_0: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_0 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_0 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1);
DATAPATH_1: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_2 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_3 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_2 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_3);
DATAPATH_2: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_4 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_5 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_4 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_5);
DATAPATH_3: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_6 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_7 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_6 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_7);
DATAPATH_4: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_8 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_9 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_4(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_4(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_4(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_4(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_4(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_8 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_9);
DATAPATH_5: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_10 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_11 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_5(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_5(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_5(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_5(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_5(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_10 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_11);
DATAPATH_6: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_12 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_13 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_6(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_6(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_6(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_6(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_6(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_12 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_13);
DATAPATH_7: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_14 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_15 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_7(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_7(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_7(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_7(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_7(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_14 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_15);
DATAPATH_8: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_16 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_17 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_8(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_8(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_8(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_8(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_8(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_16 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_17);
DATAPATH_9: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_18 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_19 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_9(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_9(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_9(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_9(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_9(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_18 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_19);
DATAPATH_10: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_20 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_21 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_10(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_10(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_10(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_10(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_10(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_20 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_21);
DATAPATH_11: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_22 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_23 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_11(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_11(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_11(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_11(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_11(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_22 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_23);
DATAPATH_12: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_24 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_25 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_12(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_12(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_12(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_12(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_12(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_24 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_25);
DATAPATH_13: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_26 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_27 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_13(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_13(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_13(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_13(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_13(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_26 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_27);
DATAPATH_14: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_28 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_29 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_14(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_14(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_14(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_14(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_14(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_28 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_29);
DATAPATH_15: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_30 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_31 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_15(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_15(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_15(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_15(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_15(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_30 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_31);
DATAPATH_16: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_32 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_33 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_16(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_16(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_16(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_16(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_16(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_32 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_33);
DATAPATH_17: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_34 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_35 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_17(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_17(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_17(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_17(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_17(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_34 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_35);
DATAPATH_18: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_36 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_37 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_18(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_18(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_18(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_18(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_18(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_36 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_37);
DATAPATH_19: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_38 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_39 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_19(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_19(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_19(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_19(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_19(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_38 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_39);
DATAPATH_20: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_40 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_41 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_20(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_20(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_20(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_20(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_20(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_40 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_41);
DATAPATH_21: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_42 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_43 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_21(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_21(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_21(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_21(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_21(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_42 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_43);
DATAPATH_22: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_44 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_45 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_22(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_22(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_22(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_22(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_22(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_44 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_45);
DATAPATH_23: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_46 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_47 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_23(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_23(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_23(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_23(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_23(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_46 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_47);
DATAPATH_24: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_48 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_49 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_24(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_24(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_24(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_24(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_24(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_48 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_49);
DATAPATH_25: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_50 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_51 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_25(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_25(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_25(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_25(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_25(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_50 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_51);
DATAPATH_26: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_52 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_53 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_26(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_26(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_26(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_26(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_26(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_52 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_53);
DATAPATH_27: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_54 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_55 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_27(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_27(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_27(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_27(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_27(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_54 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_55);
DATAPATH_28: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_56 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_57 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_28(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_28(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_28(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_28(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_28(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_56 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_57);
DATAPATH_29: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_58 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_59 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_29(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_29(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_29(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_29(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_29(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_58 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_59);
DATAPATH_30: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_60 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_61 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_30(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_30(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_30(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_30(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_30(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_60 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_61);
DATAPATH_31: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_62 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_63 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_31(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_31(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_31(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_31(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_31(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_62 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_63);
DATAPATH_32: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_64 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_65 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_32(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_32(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_32(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_32(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_32(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_64 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_65);
DATAPATH_33: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_66 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_67 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_33(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_33(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_33(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_33(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_33(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_66 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_67);
DATAPATH_34: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_68 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_69 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_34(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_34(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_34(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_34(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_34(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_68 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_69);
DATAPATH_35: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_70 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_71 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_35(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_35(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_35(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_35(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_35(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_70 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_71);
DATAPATH_36: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_72 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_73 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_36(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_36(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_36(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_36(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_36(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_72 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_73);
DATAPATH_37: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_74 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_75 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_37(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_37(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_37(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_37(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_37(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_74 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_75);
DATAPATH_38: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_76 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_77 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_38(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_38(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_38(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_38(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_38(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_76 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_77);
DATAPATH_39: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_78 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_79 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_39(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_39(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_39(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_39(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_39(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_78 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_79);
DATAPATH_40: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_80 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_81 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_40(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_40(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_40(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_40(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_40(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_80 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_81);
DATAPATH_41: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_82 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_83 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_41(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_41(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_41(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_41(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_41(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_82 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_83);
DATAPATH_42: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_84 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_85 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_42(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_42(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_42(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_42(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_42(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_84 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_85);
DATAPATH_43: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_86 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_87 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_43(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_43(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_43(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_43(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_43(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_86 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_87);
DATAPATH_44: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_88 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_89 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_44(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_44(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_44(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_44(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_44(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_88 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_89);
DATAPATH_45: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_90 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_91 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_45(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_45(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_45(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_45(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_45(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_90 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_91);
DATAPATH_46: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_92 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_93 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_46(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_46(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_46(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_46(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_46(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_92 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_93);
DATAPATH_47: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_94 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_95 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_47(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_47(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_47(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_47(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_47(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_94 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_95);
DATAPATH_48: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_96 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_97 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_48(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_48(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_48(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_48(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_48(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_96 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_97);
DATAPATH_49: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_98 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_99 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_49(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_49(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_49(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_49(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_49(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_98 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_99);
DATAPATH_50: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_100 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_101 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_50(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_50(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_50(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_50(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_50(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_100 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_101);
DATAPATH_51: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_102 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_103 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_51(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_51(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_51(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_51(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_51(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_102 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_103);
DATAPATH_52: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_104 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_105 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_52(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_52(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_52(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_52(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_52(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_104 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_105);
DATAPATH_53: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_106 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_107 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_53(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_53(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_53(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_53(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_53(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_106 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_107);
DATAPATH_54: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_108 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_109 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_54(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_54(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_54(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_54(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_54(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_108 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_109);
DATAPATH_55: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_110 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_111 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_55(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_55(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_55(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_55(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_55(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_110 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_111);
DATAPATH_56: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_112 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_113 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_56(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_56(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_56(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_56(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_56(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_112 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_113);
DATAPATH_57: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_114 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_115 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_57(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_57(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_57(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_57(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_57(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_114 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_115);
DATAPATH_58: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_116 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_117 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_58(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_58(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_58(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_58(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_58(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_116 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_117);
DATAPATH_59: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_118 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_119 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_59(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_59(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_59(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_59(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_59(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_118 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_119);
DATAPATH_60: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_120 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_121 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_60(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_60(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_60(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_60(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_60(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_120 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_121);
DATAPATH_61: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_122 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_123 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_61(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_61(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_61(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_61(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_61(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_122 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_123);
DATAPATH_62: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_124 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_125 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_62(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_62(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_62(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_62(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_62(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_124 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_125);
DATAPATH_63: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_126 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_127 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_63(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_63(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_63(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_63(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_63(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_126 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_127);
DATAPATH_64: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_128 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_129 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_64(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_64(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_64(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_64(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_64(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_128 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_129);
DATAPATH_65: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_130 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_131 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_65(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_65(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_65(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_65(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_65(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_130 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_131);
DATAPATH_66: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_132 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_133 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_66(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_66(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_66(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_66(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_66(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_132 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_133);
DATAPATH_67: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_134 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_135 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_67(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_67(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_67(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_67(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_67(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_134 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_135);
DATAPATH_68: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_136 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_137 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_68(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_68(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_68(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_68(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_68(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_136 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_137);
DATAPATH_69: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_138 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_139 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_69(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_69(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_69(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_69(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_69(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_138 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_139);
DATAPATH_70: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_140 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_141 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_70(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_70(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_70(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_70(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_70(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_140 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_141);
DATAPATH_71: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_142 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_143 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_71(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_71(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_71(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_71(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_71(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_142 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_143);
DATAPATH_72: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_144 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_145 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_72(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_72(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_72(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_72(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_72(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_144 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_145);
DATAPATH_73: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_146 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_147 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_73(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_73(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_73(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_73(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_73(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_146 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_147);
DATAPATH_74: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_148 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_149 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_74(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_74(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_74(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_74(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_74(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_148 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_149);
DATAPATH_75: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_150 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_151 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_75(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_75(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_75(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_75(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_75(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_150 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_151);
DATAPATH_76: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_152 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_153 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_76(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_76(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_76(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_76(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_76(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_152 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_153);
DATAPATH_77: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_154 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_155 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_77(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_77(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_77(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_77(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_77(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_154 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_155);
DATAPATH_78: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_156 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_157 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_78(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_78(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_78(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_78(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_78(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_156 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_157);
DATAPATH_79: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_158 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_159 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_79(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_79(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_79(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_79(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_79(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_158 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_159);
DATAPATH_80: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_160 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_161 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_80(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_80(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_80(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_80(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_80(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_160 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_161);
DATAPATH_81: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_162 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_163 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_81(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_81(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_81(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_81(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_81(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_162 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_163);
DATAPATH_82: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_164 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_165 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_82(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_82(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_82(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_82(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_82(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_164 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_165);
DATAPATH_83: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_166 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_167 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_83(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_83(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_83(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_83(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_83(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_166 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_167);
DATAPATH_84: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_168 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_169 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_84(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_84(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_84(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_84(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_84(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_168 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_169);
DATAPATH_85: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_170 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_171 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_85(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_85(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_85(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_85(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_85(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_170 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_171);
DATAPATH_86: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_172 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_173 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_86(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_86(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_86(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_86(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_86(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_172 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_173);
DATAPATH_87: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_174 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_175 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_87(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_87(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_87(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_87(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_87(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_174 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_175);
DATAPATH_88: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_176 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_177 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_88(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_88(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_88(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_88(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_88(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_176 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_177);
DATAPATH_89: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_178 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_179 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_89(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_89(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_89(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_89(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_89(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_178 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_179);
DATAPATH_90: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_180 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_181 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_90(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_90(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_90(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_90(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_90(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_180 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_181);
DATAPATH_91: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_182 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_183 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_91(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_91(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_91(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_91(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_91(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_182 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_183);
DATAPATH_92: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_184 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_185 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_92(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_92(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_92(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_92(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_92(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_184 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_185);
DATAPATH_93: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_186 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_187 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_93(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_93(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_93(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_93(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_93(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_186 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_187);
DATAPATH_94: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_188 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_189 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_94(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_94(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_94(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_94(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_94(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_188 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_189);
DATAPATH_95: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_190 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_191 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_95(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_95(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_95(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_95(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_95(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_190 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_191);
DATAPATH_96: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_192 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_193 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_96(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_96(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_96(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_96(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_96(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_192 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_193);
DATAPATH_97: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_194 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_195 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_97(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_97(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_97(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_97(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_97(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_194 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_195);
DATAPATH_98: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_196 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_197 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_98(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_98(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_98(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_98(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_98(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_196 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_197);
DATAPATH_99: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_198 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_199 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_99(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_99(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_99(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_99(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_99(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_198 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_199);
DATAPATH_100: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_200 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_201 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_100(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_100(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_100(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_100(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_100(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_200 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_201);
DATAPATH_101: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_202 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_203 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_101(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_101(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_101(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_101(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_101(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_202 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_203);
DATAPATH_102: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_204 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_205 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_102(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_102(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_102(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_102(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_102(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_204 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_205);
DATAPATH_103: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_206 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_207 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_103(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_103(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_103(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_103(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_103(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_206 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_207);
DATAPATH_104: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_208 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_209 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_104(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_104(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_104(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_104(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_104(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_208 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_209);
DATAPATH_105: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_210 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_211 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_105(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_105(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_105(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_105(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_105(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_210 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_211);
DATAPATH_106: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_212 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_213 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_106(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_106(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_106(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_106(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_106(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_212 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_213);
DATAPATH_107: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_214 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_215 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_107(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_107(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_107(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_107(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_107(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_214 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_215);
DATAPATH_108: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_216 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_217 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_108(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_108(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_108(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_108(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_108(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_216 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_217);
DATAPATH_109: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_218 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_219 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_109(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_109(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_109(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_109(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_109(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_218 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_219);
DATAPATH_110: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_220 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_221 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_110(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_110(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_110(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_110(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_110(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_220 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_221);
DATAPATH_111: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_222 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_223 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_111(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_111(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_111(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_111(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_111(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_222 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_223);
DATAPATH_112: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_224 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_225 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_112(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_112(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_112(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_112(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_112(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_224 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_225);
DATAPATH_113: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_226 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_227 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_113(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_113(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_113(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_113(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_113(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_226 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_227);
DATAPATH_114: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_228 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_229 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_114(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_114(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_114(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_114(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_114(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_228 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_229);
DATAPATH_115: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_230 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_231 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_115(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_115(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_115(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_115(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_115(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_230 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_231);
DATAPATH_116: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_232 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_233 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_116(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_116(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_116(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_116(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_116(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_232 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_233);
DATAPATH_117: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_234 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_235 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_117(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_117(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_117(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_117(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_117(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_234 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_235);
DATAPATH_118: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_236 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_237 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_118(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_118(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_118(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_118(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_118(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_236 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_237);
DATAPATH_119: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_238 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_239 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_119(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_119(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_119(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_119(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_119(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_238 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_239);
DATAPATH_120: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_240 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_241 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_120(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_120(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_120(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_120(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_120(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_240 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_241);
DATAPATH_121: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_242 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_243 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_121(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_121(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_121(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_121(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_121(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_242 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_243);
DATAPATH_122: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_244 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_245 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_122(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_122(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_122(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_122(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_122(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_244 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_245);
DATAPATH_123: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_246 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_247 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_123(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_123(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_123(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_123(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_123(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_246 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_247);
DATAPATH_124: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_248 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_249 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_124(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_124(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_124(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_124(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_124(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_248 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_249);
DATAPATH_125: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_250 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_251 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_125(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_125(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_125(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_125(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_125(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_250 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_251);
DATAPATH_126: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_252 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_253 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_126(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_126(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_126(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_126(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_126(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_252 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_253);
DATAPATH_127: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_254 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_255 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_127(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_127(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_127(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_127(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_127(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_254 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_255);
DATAPATH_128: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_256 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_257 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_128(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_128(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_128(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_128(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_128(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_256 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_257);
DATAPATH_129: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_258 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_259 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_129(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_129(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_129(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_129(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_129(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_258 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_259);
DATAPATH_130: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_260 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_261 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_130(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_130(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_130(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_130(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_130(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_260 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_261);
DATAPATH_131: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_262 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_263 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_131(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_131(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_131(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_131(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_131(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_262 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_263);
DATAPATH_132: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_264 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_265 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_132(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_132(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_132(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_132(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_132(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_264 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_265);
DATAPATH_133: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_266 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_267 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_133(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_133(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_133(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_133(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_133(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_266 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_267);
DATAPATH_134: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_268 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_269 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_134(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_134(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_134(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_134(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_134(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_268 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_269);
DATAPATH_135: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_270 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_271 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_135(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_135(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_135(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_135(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_135(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_270 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_271);
DATAPATH_136: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_272 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_273 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_136(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_136(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_136(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_136(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_136(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_272 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_273);
DATAPATH_137: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_274 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_275 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_137(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_137(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_137(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_137(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_137(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_274 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_275);
DATAPATH_138: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_276 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_277 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_138(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_138(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_138(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_138(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_138(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_276 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_277);
DATAPATH_139: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_278 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_279 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_139(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_139(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_139(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_139(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_139(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_278 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_279);
DATAPATH_140: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_280 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_281 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_140(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_140(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_140(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_140(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_140(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_280 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_281);
DATAPATH_141: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_282 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_283 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_141(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_141(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_141(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_141(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_141(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_282 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_283);
DATAPATH_142: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_284 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_285 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_142(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_142(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_142(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_142(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_142(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_284 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_285);
DATAPATH_143: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_286 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_287 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_143(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_143(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_143(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_143(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_143(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_286 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_287);
DATAPATH_144: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_288 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_289 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_144(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_144(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_144(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_144(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_144(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_288 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_289);
DATAPATH_145: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_290 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_291 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_145(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_145(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_145(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_145(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_145(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_290 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_291);
DATAPATH_146: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_292 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_293 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_146(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_146(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_146(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_146(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_146(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_292 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_293);
DATAPATH_147: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_294 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_295 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_147(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_147(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_147(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_147(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_147(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_294 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_295);
DATAPATH_148: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_296 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_297 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_148(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_148(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_148(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_148(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_148(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_296 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_297);
DATAPATH_149: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_298 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_299 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_149(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_149(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_149(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_149(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_149(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_298 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_299);
DATAPATH_150: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_300 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_301 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_150(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_150(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_150(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_150(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_150(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_300 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_301);
DATAPATH_151: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_302 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_303 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_151(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_151(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_151(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_151(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_151(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_302 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_303);
DATAPATH_152: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_304 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_305 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_152(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_152(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_152(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_152(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_152(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_304 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_305);
DATAPATH_153: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_306 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_307 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_153(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_153(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_153(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_153(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_153(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_306 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_307);
DATAPATH_154: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_308 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_309 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_154(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_154(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_154(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_154(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_154(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_308 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_309);
DATAPATH_155: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_310 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_311 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_155(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_155(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_155(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_155(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_155(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_310 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_311);
DATAPATH_156: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_312 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_313 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_156(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_156(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_156(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_156(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_156(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_312 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_313);
DATAPATH_157: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_314 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_315 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_157(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_157(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_157(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_157(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_157(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_314 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_315);
DATAPATH_158: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_316 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_317 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_158(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_158(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_158(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_158(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_158(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_316 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_317);
DATAPATH_159: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_318 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_319 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_159(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_159(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_159(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_159(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_159(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_318 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_319);
DATAPATH_160: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_320 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_321 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_160(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_160(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_160(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_160(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_160(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_320 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_321);
DATAPATH_161: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_322 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_323 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_161(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_161(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_161(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_161(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_161(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_322 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_323);
DATAPATH_162: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_324 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_325 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_162(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_162(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_162(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_162(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_162(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_324 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_325);
DATAPATH_163: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_326 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_327 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_163(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_163(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_163(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_163(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_163(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_326 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_327);
DATAPATH_164: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_328 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_329 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_164(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_164(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_164(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_164(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_164(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_328 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_329);
DATAPATH_165: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_330 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_331 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_165(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_165(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_165(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_165(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_165(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_330 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_331);
DATAPATH_166: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_332 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_333 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_166(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_166(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_166(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_166(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_166(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_332 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_333);
DATAPATH_167: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_334 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_335 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_167(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_167(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_167(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_167(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_167(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_334 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_335);
DATAPATH_168: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_336 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_337 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_168(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_168(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_168(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_168(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_168(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_336 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_337);
DATAPATH_169: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_338 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_339 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_169(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_169(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_169(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_169(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_169(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_338 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_339);
DATAPATH_170: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_340 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_341 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_170(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_170(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_170(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_170(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_170(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_340 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_341);
DATAPATH_171: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_342 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_343 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_171(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_171(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_171(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_171(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_171(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_342 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_343);
DATAPATH_172: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_344 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_345 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_172(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_172(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_172(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_172(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_172(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_344 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_345);
DATAPATH_173: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_346 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_347 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_173(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_173(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_173(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_173(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_173(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_346 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_347);
DATAPATH_174: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_348 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_349 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_174(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_174(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_174(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_174(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_174(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_348 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_349);
DATAPATH_175: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_350 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_351 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_175(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_175(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_175(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_175(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_175(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_350 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_351);
DATAPATH_176: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_352 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_353 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_176(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_176(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_176(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_176(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_176(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_352 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_353);
DATAPATH_177: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_354 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_355 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_177(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_177(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_177(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_177(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_177(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_354 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_355);
DATAPATH_178: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_356 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_357 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_178(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_178(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_178(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_178(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_178(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_356 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_357);
DATAPATH_179: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_358 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_359 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_179(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_179(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_179(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_179(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_179(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_358 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_359);
DATAPATH_180: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_360 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_361 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_180(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_180(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_180(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_180(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_180(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_360 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_361);
DATAPATH_181: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_362 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_363 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_181(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_181(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_181(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_181(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_181(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_362 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_363);
DATAPATH_182: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_364 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_365 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_182(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_182(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_182(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_182(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_182(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_364 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_365);
DATAPATH_183: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_366 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_367 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_183(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_183(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_183(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_183(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_183(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_366 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_367);
DATAPATH_184: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_368 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_369 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_184(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_184(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_184(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_184(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_184(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_368 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_369);
DATAPATH_185: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_370 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_371 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_185(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_185(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_185(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_185(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_185(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_370 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_371);
DATAPATH_186: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_372 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_373 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_186(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_186(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_186(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_186(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_186(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_372 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_373);
DATAPATH_187: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_374 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_375 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_187(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_187(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_187(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_187(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_187(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_374 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_375);
DATAPATH_188: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_376 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_377 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_188(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_188(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_188(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_188(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_188(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_376 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_377);
DATAPATH_189: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_378 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_379 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_189(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_189(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_189(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_189(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_189(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_378 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_379);
DATAPATH_190: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_380 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_381 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_190(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_190(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_190(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_190(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_190(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_380 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_381);
DATAPATH_191: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_382 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_383 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_191(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_191(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_191(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_191(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_191(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_382 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_383);
DATAPATH_192: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_384 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_385 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_192(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_192(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_192(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_192(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_192(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_384 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_385);
DATAPATH_193: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_386 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_387 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_193(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_193(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_193(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_193(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_193(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_386 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_387);
DATAPATH_194: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_388 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_389 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_194(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_194(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_194(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_194(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_194(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_388 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_389);
DATAPATH_195: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_390 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_391 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_195(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_195(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_195(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_195(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_195(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_390 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_391);
DATAPATH_196: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_392 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_393 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_196(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_196(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_196(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_196(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_196(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_392 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_393);
DATAPATH_197: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_394 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_395 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_197(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_197(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_197(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_197(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_197(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_394 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_395);
DATAPATH_198: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_396 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_397 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_198(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_198(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_198(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_198(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_198(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_396 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_397);
DATAPATH_199: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_398 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_399 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_199(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_199(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_199(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_199(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_199(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_398 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_399);
DATAPATH_200: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_400 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_401 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_200(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_200(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_200(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_200(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_200(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_400 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_401);
DATAPATH_201: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_402 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_403 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_201(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_201(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_201(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_201(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_201(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_402 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_403);
DATAPATH_202: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_404 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_405 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_202(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_202(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_202(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_202(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_202(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_404 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_405);
DATAPATH_203: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_406 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_407 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_203(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_203(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_203(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_203(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_203(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_406 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_407);
DATAPATH_204: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_408 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_409 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_204(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_204(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_204(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_204(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_204(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_408 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_409);
DATAPATH_205: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_410 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_411 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_205(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_205(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_205(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_205(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_205(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_410 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_411);
DATAPATH_206: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_412 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_413 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_206(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_206(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_206(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_206(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_206(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_412 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_413);
DATAPATH_207: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_414 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_415 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_207(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_207(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_207(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_207(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_207(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_414 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_415);
DATAPATH_208: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_416 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_417 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_208(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_208(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_208(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_208(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_208(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_416 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_417);
DATAPATH_209: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_418 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_419 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_209(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_209(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_209(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_209(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_209(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_418 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_419);
DATAPATH_210: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_420 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_421 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_210(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_210(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_210(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_210(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_210(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_420 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_421);
DATAPATH_211: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_422 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_423 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_211(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_211(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_211(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_211(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_211(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_422 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_423);
DATAPATH_212: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_424 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_425 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_212(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_212(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_212(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_212(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_212(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_424 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_425);
DATAPATH_213: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_426 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_427 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_213(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_213(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_213(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_213(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_213(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_426 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_427);
DATAPATH_214: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_428 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_429 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_214(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_214(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_214(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_214(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_214(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_428 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_429);
DATAPATH_215: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_430 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_431 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_215(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_215(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_215(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_215(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_215(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_430 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_431);
DATAPATH_216: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_432 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_433 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_216(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_216(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_216(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_216(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_216(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_432 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_433);
DATAPATH_217: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_434 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_435 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_217(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_217(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_217(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_217(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_217(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_434 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_435);
DATAPATH_218: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_436 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_437 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_218(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_218(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_218(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_218(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_218(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_436 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_437);
DATAPATH_219: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_438 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_439 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_219(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_219(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_219(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_219(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_219(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_438 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_439);
DATAPATH_220: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_440 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_441 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_220(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_220(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_220(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_220(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_220(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_440 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_441);
DATAPATH_221: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_442 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_443 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_221(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_221(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_221(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_221(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_221(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_442 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_443);
DATAPATH_222: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_444 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_445 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_222(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_222(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_222(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_222(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_222(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_444 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_445);
DATAPATH_223: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_446 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_447 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_223(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_223(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_223(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_223(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_223(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_446 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_447);
DATAPATH_224: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_448 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_449 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_224(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_224(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_224(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_224(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_224(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_448 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_449);
DATAPATH_225: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_450 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_451 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_225(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_225(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_225(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_225(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_225(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_450 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_451);
DATAPATH_226: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_452 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_453 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_226(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_226(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_226(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_226(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_226(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_452 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_453);
DATAPATH_227: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_454 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_455 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_227(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_227(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_227(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_227(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_227(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_454 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_455);
DATAPATH_228: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_456 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_457 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_228(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_228(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_228(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_228(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_228(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_456 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_457);
DATAPATH_229: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_458 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_459 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_229(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_229(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_229(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_229(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_229(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_458 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_459);
DATAPATH_230: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_460 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_461 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_230(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_230(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_230(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_230(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_230(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_460 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_461);
DATAPATH_231: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_462 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_463 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_231(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_231(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_231(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_231(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_231(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_462 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_463);
DATAPATH_232: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_464 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_465 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_232(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_232(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_232(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_232(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_232(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_464 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_465);
DATAPATH_233: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_466 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_467 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_233(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_233(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_233(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_233(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_233(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_466 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_467);
DATAPATH_234: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_468 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_469 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_234(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_234(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_234(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_234(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_234(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_468 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_469);
DATAPATH_235: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_470 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_471 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_235(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_235(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_235(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_235(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_235(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_470 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_471);
DATAPATH_236: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_472 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_473 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_236(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_236(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_236(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_236(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_236(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_472 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_473);
DATAPATH_237: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_474 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_475 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_237(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_237(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_237(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_237(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_237(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_474 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_475);
DATAPATH_238: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_476 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_477 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_238(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_238(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_238(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_238(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_238(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_476 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_477);
DATAPATH_239: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_478 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_479 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_239(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_239(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_239(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_239(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_239(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_478 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_479);
DATAPATH_240: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_480 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_481 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_240(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_240(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_240(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_240(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_240(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_480 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_481);
DATAPATH_241: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_482 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_483 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_241(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_241(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_241(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_241(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_241(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_482 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_483);
DATAPATH_242: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_484 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_485 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_242(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_242(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_242(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_242(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_242(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_484 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_485);
DATAPATH_243: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_486 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_487 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_243(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_243(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_243(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_243(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_243(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_486 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_487);
DATAPATH_244: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_488 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_489 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_244(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_244(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_244(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_244(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_244(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_488 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_489);
DATAPATH_245: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_490 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_491 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_245(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_245(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_245(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_245(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_245(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_490 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_491);
DATAPATH_246: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_492 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_493 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_246(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_246(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_246(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_246(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_246(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_492 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_493);
DATAPATH_247: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_494 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_495 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_247(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_247(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_247(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_247(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_247(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_494 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_495);
DATAPATH_248: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_496 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_497 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_248(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_248(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_248(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_248(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_248(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_496 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_497);
DATAPATH_249: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_498 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_499 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_249(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_249(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_249(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_249(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_249(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_498 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_499);
DATAPATH_250: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_500 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_501 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_250(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_250(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_250(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_250(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_250(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_500 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_501);
DATAPATH_251: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_502 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_503 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_251(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_251(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_251(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_251(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_251(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_502 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_503);
DATAPATH_252: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_504 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_505 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_252(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_252(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_252(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_252(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_252(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_504 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_505);
DATAPATH_253: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_506 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_507 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_253(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_253(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_253(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_253(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_253(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_506 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_507);
DATAPATH_254: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_508 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_509 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_254(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_254(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_254(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_254(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_254(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_508 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_509);
DATAPATH_255: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_510 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_511 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_255(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_255(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_255(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_255(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_255(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_510 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_511);
DATAPATH_256: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_512 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_513 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_256(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_256(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_256(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_256(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_256(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_512 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_513);
DATAPATH_257: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_514 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_515 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_257(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_257(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_257(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_257(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_257(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_514 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_515);
DATAPATH_258: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_516 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_517 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_258(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_258(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_258(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_258(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_258(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_516 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_517);
DATAPATH_259: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_518 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_519 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_259(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_259(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_259(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_259(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_259(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_518 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_519);
DATAPATH_260: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_520 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_521 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_260(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_260(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_260(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_260(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_260(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_520 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_521);
DATAPATH_261: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_522 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_523 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_261(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_261(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_261(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_261(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_261(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_522 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_523);
DATAPATH_262: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_524 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_525 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_262(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_262(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_262(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_262(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_262(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_524 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_525);
DATAPATH_263: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_526 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_527 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_263(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_263(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_263(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_263(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_263(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_526 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_527);
DATAPATH_264: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_528 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_529 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_264(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_264(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_264(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_264(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_264(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_528 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_529);
DATAPATH_265: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_530 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_531 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_265(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_265(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_265(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_265(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_265(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_530 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_531);
DATAPATH_266: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_532 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_533 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_266(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_266(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_266(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_266(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_266(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_532 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_533);
DATAPATH_267: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_534 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_535 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_267(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_267(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_267(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_267(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_267(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_534 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_535);
DATAPATH_268: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_536 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_537 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_268(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_268(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_268(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_268(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_268(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_536 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_537);
DATAPATH_269: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_538 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_539 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_269(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_269(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_269(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_269(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_269(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_538 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_539);
DATAPATH_270: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_540 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_541 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_270(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_270(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_270(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_270(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_270(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_540 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_541);
DATAPATH_271: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_542 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_543 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_271(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_271(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_271(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_271(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_271(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_542 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_543);
DATAPATH_272: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_544 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_545 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_272(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_272(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_272(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_272(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_272(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_544 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_545);
DATAPATH_273: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_546 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_547 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_273(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_273(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_273(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_273(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_273(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_546 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_547);
DATAPATH_274: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_548 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_549 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_274(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_274(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_274(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_274(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_274(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_548 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_549);
DATAPATH_275: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_550 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_551 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_275(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_275(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_275(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_275(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_275(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_550 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_551);
DATAPATH_276: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_552 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_553 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_276(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_276(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_276(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_276(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_276(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_552 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_553);
DATAPATH_277: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_554 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_555 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_277(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_277(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_277(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_277(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_277(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_554 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_555);
DATAPATH_278: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_556 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_557 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_278(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_278(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_278(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_278(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_278(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_556 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_557);
DATAPATH_279: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_558 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_559 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_279(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_279(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_279(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_279(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_279(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_558 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_559);
DATAPATH_280: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_560 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_561 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_280(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_280(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_280(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_280(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_280(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_560 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_561);
DATAPATH_281: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_562 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_563 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_281(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_281(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_281(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_281(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_281(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_562 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_563);
DATAPATH_282: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_564 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_565 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_282(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_282(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_282(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_282(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_282(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_564 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_565);
DATAPATH_283: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_566 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_567 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_283(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_283(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_283(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_283(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_283(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_566 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_567);
DATAPATH_284: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_568 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_569 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_284(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_284(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_284(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_284(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_284(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_568 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_569);
DATAPATH_285: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_570 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_571 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_285(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_285(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_285(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_285(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_285(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_570 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_571);
DATAPATH_286: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_572 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_573 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_286(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_286(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_286(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_286(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_286(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_572 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_573);
DATAPATH_287: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_574 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_575 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_287(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_287(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_287(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_287(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_287(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_574 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_575);
DATAPATH_288: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_576 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_577 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_288(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_288(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_288(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_288(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_288(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_576 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_577);
DATAPATH_289: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_578 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_579 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_289(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_289(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_289(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_289(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_289(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_578 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_579);
DATAPATH_290: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_580 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_581 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_290(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_290(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_290(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_290(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_290(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_580 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_581);
DATAPATH_291: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_582 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_583 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_291(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_291(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_291(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_291(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_291(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_582 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_583);
DATAPATH_292: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_584 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_585 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_292(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_292(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_292(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_292(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_292(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_584 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_585);
DATAPATH_293: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_586 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_587 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_293(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_293(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_293(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_293(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_293(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_586 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_587);
DATAPATH_294: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_588 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_589 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_294(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_294(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_294(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_294(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_294(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_588 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_589);
DATAPATH_295: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_590 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_591 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_295(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_295(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_295(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_295(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_295(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_590 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_591);
DATAPATH_296: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_592 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_593 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_296(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_296(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_296(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_296(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_296(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_592 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_593);
DATAPATH_297: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_594 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_595 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_297(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_297(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_297(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_297(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_297(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_594 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_595);
DATAPATH_298: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_596 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_597 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_298(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_298(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_298(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_298(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_298(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_596 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_597);
DATAPATH_299: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_598 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_599 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_299(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_299(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_299(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_299(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_299(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_598 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_599);
DATAPATH_300: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_600 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_601 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_300(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_300(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_300(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_300(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_300(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_600 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_601);
DATAPATH_301: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_602 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_603 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_301(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_301(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_301(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_301(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_301(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_602 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_603);
DATAPATH_302: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_604 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_605 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_302(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_302(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_302(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_302(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_302(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_604 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_605);
DATAPATH_303: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_606 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_607 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_303(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_303(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_303(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_303(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_303(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_606 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_607);
DATAPATH_304: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_608 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_609 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_304(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_304(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_304(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_304(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_304(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_608 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_609);
DATAPATH_305: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_610 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_611 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_305(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_305(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_305(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_305(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_305(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_610 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_611);
DATAPATH_306: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_612 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_613 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_306(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_306(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_306(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_306(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_306(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_612 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_613);
DATAPATH_307: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_614 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_615 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_307(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_307(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_307(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_307(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_307(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_614 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_615);
DATAPATH_308: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_616 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_617 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_308(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_308(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_308(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_308(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_308(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_616 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_617);
DATAPATH_309: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_618 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_619 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_309(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_309(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_309(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_309(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_309(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_618 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_619);
DATAPATH_310: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_620 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_621 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_310(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_310(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_310(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_310(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_310(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_620 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_621);
DATAPATH_311: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_622 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_623 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_311(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_311(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_311(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_311(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_311(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_622 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_623);
DATAPATH_312: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_624 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_625 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_312(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_312(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_312(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_312(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_312(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_624 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_625);
DATAPATH_313: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_626 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_627 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_313(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_313(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_313(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_313(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_313(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_626 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_627);
DATAPATH_314: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_628 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_629 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_314(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_314(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_314(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_314(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_314(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_628 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_629);
DATAPATH_315: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_630 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_631 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_315(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_315(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_315(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_315(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_315(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_630 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_631);
DATAPATH_316: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_632 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_633 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_316(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_316(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_316(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_316(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_316(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_632 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_633);
DATAPATH_317: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_634 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_635 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_317(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_317(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_317(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_317(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_317(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_634 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_635);
DATAPATH_318: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_636 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_637 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_318(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_318(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_318(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_318(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_318(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_636 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_637);
DATAPATH_319: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_638 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_639 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_319(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_319(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_319(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_319(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_319(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_638 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_639);
DATAPATH_320: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_640 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_641 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_320(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_320(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_320(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_320(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_320(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_640 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_641);
DATAPATH_321: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_642 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_643 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_321(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_321(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_321(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_321(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_321(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_642 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_643);
DATAPATH_322: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_644 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_645 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_322(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_322(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_322(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_322(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_322(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_644 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_645);
DATAPATH_323: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_646 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_647 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_323(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_323(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_323(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_323(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_323(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_646 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_647);
DATAPATH_324: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_648 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_649 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_324(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_324(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_324(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_324(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_324(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_648 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_649);
DATAPATH_325: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_650 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_651 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_325(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_325(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_325(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_325(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_325(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_650 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_651);
DATAPATH_326: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_652 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_653 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_326(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_326(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_326(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_326(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_326(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_652 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_653);
DATAPATH_327: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_654 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_655 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_327(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_327(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_327(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_327(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_327(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_654 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_655);
DATAPATH_328: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_656 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_657 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_328(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_328(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_328(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_328(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_328(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_656 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_657);
DATAPATH_329: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_658 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_659 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_329(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_329(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_329(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_329(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_329(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_658 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_659);
DATAPATH_330: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_660 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_661 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_330(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_330(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_330(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_330(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_330(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_660 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_661);
DATAPATH_331: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_662 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_663 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_331(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_331(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_331(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_331(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_331(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_662 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_663);
DATAPATH_332: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_664 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_665 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_332(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_332(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_332(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_332(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_332(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_664 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_665);
DATAPATH_333: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_666 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_667 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_333(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_333(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_333(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_333(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_333(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_666 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_667);
DATAPATH_334: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_668 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_669 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_334(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_334(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_334(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_334(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_334(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_668 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_669);
DATAPATH_335: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_670 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_671 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_335(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_335(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_335(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_335(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_335(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_670 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_671);
DATAPATH_336: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_672 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_673 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_336(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_336(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_336(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_336(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_336(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_672 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_673);
DATAPATH_337: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_674 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_675 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_337(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_337(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_337(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_337(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_337(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_674 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_675);
DATAPATH_338: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_676 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_677 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_338(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_338(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_338(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_338(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_338(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_676 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_677);
DATAPATH_339: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_678 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_679 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_339(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_339(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_339(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_339(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_339(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_678 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_679);
DATAPATH_340: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_680 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_681 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_340(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_340(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_340(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_340(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_340(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_680 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_681);
DATAPATH_341: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_682 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_683 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_341(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_341(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_341(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_341(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_341(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_682 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_683);
DATAPATH_342: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_684 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_685 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_342(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_342(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_342(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_342(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_342(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_684 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_685);
DATAPATH_343: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_686 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_687 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_343(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_343(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_343(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_343(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_343(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_686 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_687);
DATAPATH_344: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_688 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_689 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_344(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_344(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_344(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_344(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_344(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_688 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_689);
DATAPATH_345: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_690 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_691 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_345(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_345(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_345(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_345(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_345(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_690 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_691);
DATAPATH_346: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_692 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_693 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_346(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_346(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_346(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_346(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_346(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_692 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_693);
DATAPATH_347: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_694 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_695 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_347(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_347(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_347(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_347(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_347(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_694 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_695);
DATAPATH_348: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_696 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_697 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_348(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_348(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_348(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_348(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_348(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_696 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_697);
DATAPATH_349: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_698 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_699 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_349(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_349(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_349(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_349(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_349(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_698 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_699);
DATAPATH_350: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_700 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_701 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_350(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_350(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_350(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_350(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_350(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_700 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_701);
DATAPATH_351: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_702 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_703 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_351(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_351(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_351(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_351(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_351(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_702 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_703);
DATAPATH_352: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_704 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_705 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_352(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_352(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_352(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_352(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_352(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_704 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_705);
DATAPATH_353: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_706 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_707 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_353(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_353(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_353(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_353(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_353(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_706 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_707);
DATAPATH_354: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_708 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_709 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_354(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_354(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_354(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_354(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_354(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_708 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_709);
DATAPATH_355: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_710 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_711 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_355(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_355(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_355(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_355(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_355(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_710 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_711);
DATAPATH_356: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_712 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_713 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_356(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_356(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_356(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_356(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_356(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_712 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_713);
DATAPATH_357: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_714 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_715 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_357(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_357(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_357(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_357(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_357(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_714 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_715);
DATAPATH_358: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_716 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_717 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_358(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_358(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_358(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_358(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_358(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_716 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_717);
DATAPATH_359: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_718 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_719 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_359(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_359(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_359(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_359(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_359(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_718 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_719);
DATAPATH_360: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_720 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_721 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_360(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_360(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_360(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_360(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_360(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_720 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_721);
DATAPATH_361: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_722 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_723 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_361(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_361(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_361(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_361(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_361(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_722 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_723);
DATAPATH_362: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_724 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_725 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_362(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_362(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_362(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_362(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_362(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_724 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_725);
DATAPATH_363: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_726 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_727 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_363(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_363(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_363(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_363(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_363(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_726 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_727);
DATAPATH_364: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_728 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_729 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_364(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_364(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_364(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_364(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_364(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_728 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_729);
DATAPATH_365: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_730 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_731 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_365(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_365(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_365(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_365(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_365(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_730 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_731);
DATAPATH_366: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_732 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_733 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_366(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_366(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_366(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_366(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_366(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_732 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_733);
DATAPATH_367: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_734 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_735 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_367(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_367(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_367(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_367(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_367(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_734 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_735);
DATAPATH_368: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_736 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_737 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_368(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_368(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_368(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_368(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_368(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_736 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_737);
DATAPATH_369: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_738 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_739 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_369(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_369(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_369(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_369(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_369(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_738 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_739);
DATAPATH_370: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_740 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_741 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_370(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_370(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_370(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_370(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_370(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_740 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_741);
DATAPATH_371: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_742 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_743 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_371(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_371(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_371(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_371(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_371(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_742 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_743);
DATAPATH_372: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_744 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_745 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_372(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_372(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_372(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_372(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_372(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_744 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_745);
DATAPATH_373: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_746 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_747 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_373(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_373(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_373(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_373(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_373(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_746 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_747);
DATAPATH_374: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_748 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_749 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_374(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_374(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_374(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_374(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_374(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_748 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_749);
DATAPATH_375: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_750 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_751 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_375(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_375(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_375(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_375(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_375(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_750 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_751);
DATAPATH_376: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_752 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_753 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_376(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_376(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_376(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_376(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_376(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_752 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_753);
DATAPATH_377: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_754 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_755 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_377(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_377(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_377(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_377(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_377(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_754 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_755);
DATAPATH_378: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_756 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_757 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_378(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_378(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_378(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_378(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_378(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_756 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_757);
DATAPATH_379: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_758 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_759 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_379(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_379(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_379(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_379(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_379(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_758 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_759);
DATAPATH_380: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_760 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_761 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_380(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_380(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_380(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_380(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_380(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_760 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_761);
DATAPATH_381: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_762 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_763 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_381(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_381(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_381(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_381(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_381(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_762 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_763);
DATAPATH_382: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_764 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_765 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_382(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_382(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_382(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_382(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_382(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_764 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_765);
DATAPATH_383: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_766 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_767 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_383(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_383(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_383(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_383(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_383(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_766 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_767);
DATAPATH_384: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_768 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_769 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_384(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_384(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_384(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_384(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_384(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_768 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_769);
DATAPATH_385: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_770 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_771 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_385(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_385(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_385(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_385(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_385(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_770 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_771);
DATAPATH_386: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_772 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_773 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_386(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_386(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_386(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_386(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_386(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_772 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_773);
DATAPATH_387: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_774 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_775 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_387(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_387(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_387(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_387(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_387(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_774 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_775);
DATAPATH_388: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_776 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_777 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_388(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_388(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_388(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_388(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_388(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_776 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_777);
DATAPATH_389: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_778 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_779 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_389(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_389(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_389(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_389(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_389(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_778 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_779);
DATAPATH_390: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_780 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_781 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_390(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_390(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_390(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_390(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_390(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_780 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_781);
DATAPATH_391: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_782 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_783 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_391(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_391(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_391(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_391(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_391(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_782 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_783);
DATAPATH_392: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_784 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_785 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_392(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_392(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_392(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_392(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_392(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_784 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_785);
DATAPATH_393: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_786 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_787 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_393(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_393(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_393(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_393(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_393(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_786 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_787);
DATAPATH_394: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_788 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_789 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_394(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_394(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_394(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_394(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_394(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_788 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_789);
DATAPATH_395: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_790 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_791 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_395(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_395(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_395(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_395(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_395(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_790 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_791);
DATAPATH_396: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_792 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_793 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_396(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_396(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_396(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_396(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_396(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_792 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_793);
DATAPATH_397: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_794 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_795 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_397(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_397(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_397(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_397(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_397(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_794 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_795);
DATAPATH_398: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_796 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_797 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_398(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_398(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_398(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_398(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_398(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_796 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_797);
DATAPATH_399: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_798 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_799 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_399(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_399(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_399(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_399(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_399(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_798 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_799);
DATAPATH_400: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_800 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_801 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_400(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_400(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_400(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_400(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_400(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_800 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_801);
DATAPATH_401: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_802 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_803 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_401(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_401(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_401(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_401(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_401(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_802 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_803);
DATAPATH_402: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_804 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_805 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_402(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_402(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_402(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_402(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_402(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_804 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_805);
DATAPATH_403: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_806 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_807 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_403(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_403(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_403(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_403(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_403(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_806 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_807);
DATAPATH_404: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_808 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_809 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_404(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_404(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_404(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_404(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_404(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_808 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_809);
DATAPATH_405: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_810 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_811 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_405(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_405(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_405(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_405(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_405(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_810 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_811);
DATAPATH_406: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_812 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_813 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_406(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_406(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_406(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_406(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_406(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_812 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_813);
DATAPATH_407: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_814 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_815 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_407(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_407(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_407(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_407(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_407(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_814 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_815);
DATAPATH_408: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_816 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_817 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_408(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_408(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_408(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_408(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_408(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_816 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_817);
DATAPATH_409: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_818 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_819 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_409(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_409(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_409(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_409(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_409(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_818 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_819);
DATAPATH_410: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_820 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_821 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_410(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_410(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_410(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_410(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_410(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_820 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_821);
DATAPATH_411: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_822 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_823 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_411(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_411(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_411(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_411(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_411(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_822 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_823);
DATAPATH_412: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_824 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_825 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_412(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_412(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_412(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_412(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_412(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_824 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_825);
DATAPATH_413: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_826 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_827 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_413(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_413(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_413(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_413(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_413(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_826 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_827);
DATAPATH_414: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_828 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_829 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_414(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_414(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_414(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_414(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_414(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_828 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_829);
DATAPATH_415: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_830 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_831 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_415(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_415(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_415(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_415(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_415(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_830 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_831);
DATAPATH_416: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_832 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_833 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_416(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_416(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_416(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_416(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_416(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_832 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_833);
DATAPATH_417: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_834 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_835 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_417(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_417(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_417(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_417(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_417(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_834 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_835);
DATAPATH_418: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_836 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_837 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_418(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_418(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_418(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_418(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_418(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_836 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_837);
DATAPATH_419: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_838 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_839 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_419(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_419(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_419(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_419(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_419(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_838 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_839);
DATAPATH_420: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_840 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_841 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_420(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_420(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_420(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_420(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_420(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_840 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_841);
DATAPATH_421: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_842 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_843 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_421(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_421(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_421(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_421(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_421(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_842 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_843);
DATAPATH_422: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_844 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_845 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_422(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_422(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_422(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_422(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_422(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_844 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_845);
DATAPATH_423: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_846 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_847 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_423(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_423(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_423(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_423(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_423(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_846 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_847);
DATAPATH_424: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_848 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_849 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_424(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_424(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_424(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_424(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_424(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_848 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_849);
DATAPATH_425: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_850 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_851 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_425(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_425(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_425(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_425(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_425(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_850 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_851);
DATAPATH_426: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_852 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_853 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_426(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_426(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_426(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_426(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_426(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_852 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_853);
DATAPATH_427: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_854 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_855 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_427(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_427(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_427(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_427(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_427(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_854 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_855);
DATAPATH_428: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_856 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_857 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_428(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_428(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_428(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_428(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_428(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_856 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_857);
DATAPATH_429: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_858 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_859 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_429(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_429(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_429(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_429(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_429(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_858 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_859);
DATAPATH_430: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_860 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_861 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_430(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_430(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_430(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_430(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_430(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_860 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_861);
DATAPATH_431: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_862 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_863 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_431(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_431(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_431(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_431(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_431(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_862 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_863);
DATAPATH_432: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_864 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_865 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_432(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_432(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_432(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_432(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_432(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_864 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_865);
DATAPATH_433: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_866 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_867 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_433(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_433(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_433(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_433(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_433(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_866 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_867);
DATAPATH_434: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_868 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_869 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_434(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_434(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_434(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_434(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_434(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_868 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_869);
DATAPATH_435: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_870 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_871 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_435(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_435(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_435(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_435(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_435(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_870 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_871);
DATAPATH_436: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_872 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_873 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_436(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_436(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_436(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_436(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_436(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_872 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_873);
DATAPATH_437: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_874 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_875 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_437(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_437(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_437(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_437(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_437(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_874 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_875);
DATAPATH_438: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_876 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_877 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_438(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_438(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_438(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_438(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_438(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_876 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_877);
DATAPATH_439: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_878 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_879 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_439(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_439(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_439(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_439(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_439(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_878 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_879);
DATAPATH_440: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_880 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_881 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_440(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_440(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_440(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_440(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_440(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_880 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_881);
DATAPATH_441: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_882 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_883 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_441(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_441(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_441(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_441(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_441(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_882 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_883);
DATAPATH_442: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_884 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_885 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_442(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_442(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_442(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_442(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_442(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_884 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_885);
DATAPATH_443: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_886 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_887 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_443(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_443(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_443(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_443(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_443(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_886 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_887);
DATAPATH_444: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_888 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_889 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_444(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_444(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_444(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_444(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_444(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_888 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_889);
DATAPATH_445: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_890 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_891 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_445(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_445(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_445(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_445(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_445(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_890 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_891);
DATAPATH_446: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_892 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_893 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_446(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_446(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_446(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_446(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_446(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_892 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_893);
DATAPATH_447: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_894 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_895 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_447(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_447(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_447(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_447(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_447(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_894 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_895);
DATAPATH_448: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_896 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_897 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_448(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_448(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_448(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_448(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_448(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_896 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_897);
DATAPATH_449: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_898 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_899 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_449(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_449(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_449(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_449(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_449(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_898 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_899);
DATAPATH_450: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_900 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_901 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_450(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_450(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_450(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_450(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_450(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_900 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_901);
DATAPATH_451: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_902 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_903 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_451(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_451(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_451(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_451(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_451(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_902 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_903);
DATAPATH_452: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_904 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_905 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_452(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_452(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_452(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_452(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_452(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_904 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_905);
DATAPATH_453: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_906 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_907 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_453(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_453(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_453(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_453(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_453(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_906 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_907);
DATAPATH_454: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_908 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_909 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_454(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_454(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_454(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_454(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_454(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_908 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_909);
DATAPATH_455: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_910 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_911 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_455(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_455(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_455(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_455(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_455(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_910 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_911);
DATAPATH_456: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_912 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_913 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_456(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_456(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_456(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_456(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_456(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_912 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_913);
DATAPATH_457: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_914 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_915 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_457(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_457(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_457(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_457(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_457(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_914 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_915);
DATAPATH_458: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_916 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_917 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_458(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_458(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_458(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_458(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_458(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_916 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_917);
DATAPATH_459: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_918 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_919 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_459(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_459(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_459(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_459(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_459(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_918 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_919);
DATAPATH_460: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_920 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_921 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_460(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_460(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_460(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_460(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_460(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_920 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_921);
DATAPATH_461: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_922 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_923 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_461(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_461(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_461(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_461(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_461(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_922 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_923);
DATAPATH_462: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_924 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_925 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_462(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_462(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_462(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_462(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_462(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_924 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_925);
DATAPATH_463: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_926 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_927 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_463(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_463(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_463(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_463(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_463(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_926 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_927);
DATAPATH_464: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_928 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_929 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_464(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_464(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_464(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_464(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_464(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_928 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_929);
DATAPATH_465: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_930 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_931 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_465(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_465(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_465(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_465(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_465(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_930 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_931);
DATAPATH_466: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_932 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_933 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_466(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_466(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_466(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_466(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_466(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_932 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_933);
DATAPATH_467: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_934 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_935 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_467(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_467(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_467(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_467(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_467(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_934 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_935);
DATAPATH_468: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_936 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_937 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_468(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_468(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_468(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_468(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_468(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_936 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_937);
DATAPATH_469: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_938 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_939 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_469(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_469(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_469(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_469(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_469(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_938 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_939);
DATAPATH_470: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_940 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_941 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_470(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_470(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_470(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_470(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_470(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_940 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_941);
DATAPATH_471: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_942 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_943 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_471(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_471(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_471(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_471(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_471(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_942 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_943);
DATAPATH_472: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_944 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_945 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_472(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_472(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_472(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_472(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_472(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_944 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_945);
DATAPATH_473: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_946 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_947 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_473(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_473(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_473(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_473(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_473(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_946 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_947);
DATAPATH_474: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_948 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_949 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_474(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_474(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_474(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_474(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_474(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_948 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_949);
DATAPATH_475: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_950 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_951 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_475(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_475(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_475(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_475(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_475(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_950 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_951);
DATAPATH_476: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_952 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_953 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_476(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_476(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_476(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_476(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_476(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_952 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_953);
DATAPATH_477: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_954 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_955 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_477(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_477(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_477(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_477(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_477(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_954 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_955);
DATAPATH_478: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_956 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_957 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_478(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_478(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_478(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_478(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_478(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_956 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_957);
DATAPATH_479: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_958 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_959 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_479(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_479(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_479(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_479(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_479(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_958 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_959);
DATAPATH_480: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_960 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_961 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_480(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_480(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_480(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_480(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_480(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_960 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_961);
DATAPATH_481: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_962 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_963 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_481(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_481(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_481(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_481(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_481(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_962 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_963);
DATAPATH_482: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_964 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_965 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_482(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_482(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_482(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_482(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_482(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_964 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_965);
DATAPATH_483: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_966 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_967 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_483(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_483(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_483(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_483(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_483(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_966 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_967);
DATAPATH_484: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_968 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_969 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_484(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_484(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_484(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_484(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_484(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_968 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_969);
DATAPATH_485: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_970 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_971 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_485(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_485(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_485(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_485(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_485(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_970 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_971);
DATAPATH_486: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_972 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_973 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_486(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_486(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_486(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_486(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_486(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_972 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_973);
DATAPATH_487: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_974 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_975 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_487(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_487(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_487(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_487(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_487(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_974 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_975);
DATAPATH_488: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_976 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_977 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_488(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_488(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_488(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_488(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_488(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_976 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_977);
DATAPATH_489: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_978 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_979 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_489(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_489(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_489(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_489(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_489(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_978 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_979);
DATAPATH_490: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_980 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_981 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_490(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_490(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_490(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_490(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_490(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_980 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_981);
DATAPATH_491: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_982 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_983 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_491(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_491(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_491(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_491(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_491(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_982 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_983);
DATAPATH_492: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_984 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_985 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_492(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_492(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_492(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_492(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_492(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_984 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_985);
DATAPATH_493: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_986 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_987 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_493(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_493(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_493(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_493(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_493(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_986 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_987);
DATAPATH_494: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_988 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_989 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_494(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_494(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_494(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_494(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_494(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_988 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_989);
DATAPATH_495: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_990 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_991 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_495(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_495(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_495(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_495(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_495(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_990 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_991);
DATAPATH_496: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_992 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_993 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_496(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_496(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_496(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_496(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_496(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_992 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_993);
DATAPATH_497: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_994 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_995 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_497(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_497(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_497(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_497(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_497(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_994 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_995);
DATAPATH_498: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_996 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_997 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_498(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_498(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_498(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_498(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_498(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_996 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_997);
DATAPATH_499: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_998 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_999 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_499(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_499(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_499(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_499(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_499(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_998 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_999);
DATAPATH_500: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1000 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1001 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_500(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_500(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_500(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_500(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_500(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1000 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1001);
DATAPATH_501: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1002 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1003 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_501(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_501(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_501(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_501(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_501(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1002 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1003);
DATAPATH_502: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1004 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1005 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_502(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_502(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_502(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_502(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_502(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1004 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1005);
DATAPATH_503: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1006 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1007 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_503(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_503(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_503(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_503(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_503(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1006 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1007);
DATAPATH_504: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1008 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1009 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_504(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_504(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_504(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_504(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_504(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1008 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1009);
DATAPATH_505: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1010 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1011 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_505(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_505(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_505(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_505(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_505(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1010 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1011);
DATAPATH_506: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1012 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1013 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_506(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_506(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_506(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_506(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_506(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1012 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1013);
DATAPATH_507: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1014 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1015 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_507(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_507(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_507(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_507(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_507(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1014 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1015);
DATAPATH_508: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1016 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1017 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_508(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_508(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_508(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_508(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_508(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1016 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1017);
DATAPATH_509: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1018 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1019 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_509(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_509(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_509(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_509(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_509(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1018 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1019);
DATAPATH_510: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1020 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1021 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_510(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_510(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_510(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_510(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_510(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1020 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1021);
DATAPATH_511: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_1022 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1023 ,
            DATAPATH_IN_SINE => QEP_N_10_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_10_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_511(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_511(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_511(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_511(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_511(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_10_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_10_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_1022 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1023);

UNWINDOWED_0 <= FROM_DATAPATHS_0;
UNWINDOWED_1 <= FROM_DATAPATHS_1;
UNWINDOWED_2 <= FROM_DATAPATHS_2;
UNWINDOWED_3 <= FROM_DATAPATHS_3;
UNWINDOWED_4 <= FROM_DATAPATHS_4;
UNWINDOWED_5 <= FROM_DATAPATHS_5;
UNWINDOWED_6 <= FROM_DATAPATHS_6;
UNWINDOWED_7 <= FROM_DATAPATHS_7;
UNWINDOWED_8 <= FROM_DATAPATHS_8;
UNWINDOWED_9 <= FROM_DATAPATHS_9;
UNWINDOWED_10 <= FROM_DATAPATHS_10;
UNWINDOWED_11 <= FROM_DATAPATHS_11;
UNWINDOWED_12 <= FROM_DATAPATHS_12;
UNWINDOWED_13 <= FROM_DATAPATHS_13;
UNWINDOWED_14 <= FROM_DATAPATHS_14;
UNWINDOWED_15 <= FROM_DATAPATHS_15;
UNWINDOWED_16 <= FROM_DATAPATHS_16;
UNWINDOWED_17 <= FROM_DATAPATHS_17;
UNWINDOWED_18 <= FROM_DATAPATHS_18;
UNWINDOWED_19 <= FROM_DATAPATHS_19;
UNWINDOWED_20 <= FROM_DATAPATHS_20;
UNWINDOWED_21 <= FROM_DATAPATHS_21;
UNWINDOWED_22 <= FROM_DATAPATHS_22;
UNWINDOWED_23 <= FROM_DATAPATHS_23;
UNWINDOWED_24 <= FROM_DATAPATHS_24;
UNWINDOWED_25 <= FROM_DATAPATHS_25;
UNWINDOWED_26 <= FROM_DATAPATHS_26;
UNWINDOWED_27 <= FROM_DATAPATHS_27;
UNWINDOWED_28 <= FROM_DATAPATHS_28;
UNWINDOWED_29 <= FROM_DATAPATHS_29;
UNWINDOWED_30 <= FROM_DATAPATHS_30;
UNWINDOWED_31 <= FROM_DATAPATHS_31;
UNWINDOWED_32 <= FROM_DATAPATHS_32;
UNWINDOWED_33 <= FROM_DATAPATHS_33;
UNWINDOWED_34 <= FROM_DATAPATHS_34;
UNWINDOWED_35 <= FROM_DATAPATHS_35;
UNWINDOWED_36 <= FROM_DATAPATHS_36;
UNWINDOWED_37 <= FROM_DATAPATHS_37;
UNWINDOWED_38 <= FROM_DATAPATHS_38;
UNWINDOWED_39 <= FROM_DATAPATHS_39;
UNWINDOWED_40 <= FROM_DATAPATHS_40;
UNWINDOWED_41 <= FROM_DATAPATHS_41;
UNWINDOWED_42 <= FROM_DATAPATHS_42;
UNWINDOWED_43 <= FROM_DATAPATHS_43;
UNWINDOWED_44 <= FROM_DATAPATHS_44;
UNWINDOWED_45 <= FROM_DATAPATHS_45;
UNWINDOWED_46 <= FROM_DATAPATHS_46;
UNWINDOWED_47 <= FROM_DATAPATHS_47;
UNWINDOWED_48 <= FROM_DATAPATHS_48;
UNWINDOWED_49 <= FROM_DATAPATHS_49;
UNWINDOWED_50 <= FROM_DATAPATHS_50;
UNWINDOWED_51 <= FROM_DATAPATHS_51;
UNWINDOWED_52 <= FROM_DATAPATHS_52;
UNWINDOWED_53 <= FROM_DATAPATHS_53;
UNWINDOWED_54 <= FROM_DATAPATHS_54;
UNWINDOWED_55 <= FROM_DATAPATHS_55;
UNWINDOWED_56 <= FROM_DATAPATHS_56;
UNWINDOWED_57 <= FROM_DATAPATHS_57;
UNWINDOWED_58 <= FROM_DATAPATHS_58;
UNWINDOWED_59 <= FROM_DATAPATHS_59;
UNWINDOWED_60 <= FROM_DATAPATHS_60;
UNWINDOWED_61 <= FROM_DATAPATHS_61;
UNWINDOWED_62 <= FROM_DATAPATHS_62;
UNWINDOWED_63 <= FROM_DATAPATHS_63;
UNWINDOWED_64 <= FROM_DATAPATHS_64;
UNWINDOWED_65 <= FROM_DATAPATHS_65;
UNWINDOWED_66 <= FROM_DATAPATHS_66;
UNWINDOWED_67 <= FROM_DATAPATHS_67;
UNWINDOWED_68 <= FROM_DATAPATHS_68;
UNWINDOWED_69 <= FROM_DATAPATHS_69;
UNWINDOWED_70 <= FROM_DATAPATHS_70;
UNWINDOWED_71 <= FROM_DATAPATHS_71;
UNWINDOWED_72 <= FROM_DATAPATHS_72;
UNWINDOWED_73 <= FROM_DATAPATHS_73;
UNWINDOWED_74 <= FROM_DATAPATHS_74;
UNWINDOWED_75 <= FROM_DATAPATHS_75;
UNWINDOWED_76 <= FROM_DATAPATHS_76;
UNWINDOWED_77 <= FROM_DATAPATHS_77;
UNWINDOWED_78 <= FROM_DATAPATHS_78;
UNWINDOWED_79 <= FROM_DATAPATHS_79;
UNWINDOWED_80 <= FROM_DATAPATHS_80;
UNWINDOWED_81 <= FROM_DATAPATHS_81;
UNWINDOWED_82 <= FROM_DATAPATHS_82;
UNWINDOWED_83 <= FROM_DATAPATHS_83;
UNWINDOWED_84 <= FROM_DATAPATHS_84;
UNWINDOWED_85 <= FROM_DATAPATHS_85;
UNWINDOWED_86 <= FROM_DATAPATHS_86;
UNWINDOWED_87 <= FROM_DATAPATHS_87;
UNWINDOWED_88 <= FROM_DATAPATHS_88;
UNWINDOWED_89 <= FROM_DATAPATHS_89;
UNWINDOWED_90 <= FROM_DATAPATHS_90;
UNWINDOWED_91 <= FROM_DATAPATHS_91;
UNWINDOWED_92 <= FROM_DATAPATHS_92;
UNWINDOWED_93 <= FROM_DATAPATHS_93;
UNWINDOWED_94 <= FROM_DATAPATHS_94;
UNWINDOWED_95 <= FROM_DATAPATHS_95;
UNWINDOWED_96 <= FROM_DATAPATHS_96;
UNWINDOWED_97 <= FROM_DATAPATHS_97;
UNWINDOWED_98 <= FROM_DATAPATHS_98;
UNWINDOWED_99 <= FROM_DATAPATHS_99;
UNWINDOWED_100 <= FROM_DATAPATHS_100;
UNWINDOWED_101 <= FROM_DATAPATHS_101;
UNWINDOWED_102 <= FROM_DATAPATHS_102;
UNWINDOWED_103 <= FROM_DATAPATHS_103;
UNWINDOWED_104 <= FROM_DATAPATHS_104;
UNWINDOWED_105 <= FROM_DATAPATHS_105;
UNWINDOWED_106 <= FROM_DATAPATHS_106;
UNWINDOWED_107 <= FROM_DATAPATHS_107;
UNWINDOWED_108 <= FROM_DATAPATHS_108;
UNWINDOWED_109 <= FROM_DATAPATHS_109;
UNWINDOWED_110 <= FROM_DATAPATHS_110;
UNWINDOWED_111 <= FROM_DATAPATHS_111;
UNWINDOWED_112 <= FROM_DATAPATHS_112;
UNWINDOWED_113 <= FROM_DATAPATHS_113;
UNWINDOWED_114 <= FROM_DATAPATHS_114;
UNWINDOWED_115 <= FROM_DATAPATHS_115;
UNWINDOWED_116 <= FROM_DATAPATHS_116;
UNWINDOWED_117 <= FROM_DATAPATHS_117;
UNWINDOWED_118 <= FROM_DATAPATHS_118;
UNWINDOWED_119 <= FROM_DATAPATHS_119;
UNWINDOWED_120 <= FROM_DATAPATHS_120;
UNWINDOWED_121 <= FROM_DATAPATHS_121;
UNWINDOWED_122 <= FROM_DATAPATHS_122;
UNWINDOWED_123 <= FROM_DATAPATHS_123;
UNWINDOWED_124 <= FROM_DATAPATHS_124;
UNWINDOWED_125 <= FROM_DATAPATHS_125;
UNWINDOWED_126 <= FROM_DATAPATHS_126;
UNWINDOWED_127 <= FROM_DATAPATHS_127;
UNWINDOWED_128 <= FROM_DATAPATHS_128;
UNWINDOWED_129 <= FROM_DATAPATHS_129;
UNWINDOWED_130 <= FROM_DATAPATHS_130;
UNWINDOWED_131 <= FROM_DATAPATHS_131;
UNWINDOWED_132 <= FROM_DATAPATHS_132;
UNWINDOWED_133 <= FROM_DATAPATHS_133;
UNWINDOWED_134 <= FROM_DATAPATHS_134;
UNWINDOWED_135 <= FROM_DATAPATHS_135;
UNWINDOWED_136 <= FROM_DATAPATHS_136;
UNWINDOWED_137 <= FROM_DATAPATHS_137;
UNWINDOWED_138 <= FROM_DATAPATHS_138;
UNWINDOWED_139 <= FROM_DATAPATHS_139;
UNWINDOWED_140 <= FROM_DATAPATHS_140;
UNWINDOWED_141 <= FROM_DATAPATHS_141;
UNWINDOWED_142 <= FROM_DATAPATHS_142;
UNWINDOWED_143 <= FROM_DATAPATHS_143;
UNWINDOWED_144 <= FROM_DATAPATHS_144;
UNWINDOWED_145 <= FROM_DATAPATHS_145;
UNWINDOWED_146 <= FROM_DATAPATHS_146;
UNWINDOWED_147 <= FROM_DATAPATHS_147;
UNWINDOWED_148 <= FROM_DATAPATHS_148;
UNWINDOWED_149 <= FROM_DATAPATHS_149;
UNWINDOWED_150 <= FROM_DATAPATHS_150;
UNWINDOWED_151 <= FROM_DATAPATHS_151;
UNWINDOWED_152 <= FROM_DATAPATHS_152;
UNWINDOWED_153 <= FROM_DATAPATHS_153;
UNWINDOWED_154 <= FROM_DATAPATHS_154;
UNWINDOWED_155 <= FROM_DATAPATHS_155;
UNWINDOWED_156 <= FROM_DATAPATHS_156;
UNWINDOWED_157 <= FROM_DATAPATHS_157;
UNWINDOWED_158 <= FROM_DATAPATHS_158;
UNWINDOWED_159 <= FROM_DATAPATHS_159;
UNWINDOWED_160 <= FROM_DATAPATHS_160;
UNWINDOWED_161 <= FROM_DATAPATHS_161;
UNWINDOWED_162 <= FROM_DATAPATHS_162;
UNWINDOWED_163 <= FROM_DATAPATHS_163;
UNWINDOWED_164 <= FROM_DATAPATHS_164;
UNWINDOWED_165 <= FROM_DATAPATHS_165;
UNWINDOWED_166 <= FROM_DATAPATHS_166;
UNWINDOWED_167 <= FROM_DATAPATHS_167;
UNWINDOWED_168 <= FROM_DATAPATHS_168;
UNWINDOWED_169 <= FROM_DATAPATHS_169;
UNWINDOWED_170 <= FROM_DATAPATHS_170;
UNWINDOWED_171 <= FROM_DATAPATHS_171;
UNWINDOWED_172 <= FROM_DATAPATHS_172;
UNWINDOWED_173 <= FROM_DATAPATHS_173;
UNWINDOWED_174 <= FROM_DATAPATHS_174;
UNWINDOWED_175 <= FROM_DATAPATHS_175;
UNWINDOWED_176 <= FROM_DATAPATHS_176;
UNWINDOWED_177 <= FROM_DATAPATHS_177;
UNWINDOWED_178 <= FROM_DATAPATHS_178;
UNWINDOWED_179 <= FROM_DATAPATHS_179;
UNWINDOWED_180 <= FROM_DATAPATHS_180;
UNWINDOWED_181 <= FROM_DATAPATHS_181;
UNWINDOWED_182 <= FROM_DATAPATHS_182;
UNWINDOWED_183 <= FROM_DATAPATHS_183;
UNWINDOWED_184 <= FROM_DATAPATHS_184;
UNWINDOWED_185 <= FROM_DATAPATHS_185;
UNWINDOWED_186 <= FROM_DATAPATHS_186;
UNWINDOWED_187 <= FROM_DATAPATHS_187;
UNWINDOWED_188 <= FROM_DATAPATHS_188;
UNWINDOWED_189 <= FROM_DATAPATHS_189;
UNWINDOWED_190 <= FROM_DATAPATHS_190;
UNWINDOWED_191 <= FROM_DATAPATHS_191;
UNWINDOWED_192 <= FROM_DATAPATHS_192;
UNWINDOWED_193 <= FROM_DATAPATHS_193;
UNWINDOWED_194 <= FROM_DATAPATHS_194;
UNWINDOWED_195 <= FROM_DATAPATHS_195;
UNWINDOWED_196 <= FROM_DATAPATHS_196;
UNWINDOWED_197 <= FROM_DATAPATHS_197;
UNWINDOWED_198 <= FROM_DATAPATHS_198;
UNWINDOWED_199 <= FROM_DATAPATHS_199;
UNWINDOWED_200 <= FROM_DATAPATHS_200;
UNWINDOWED_201 <= FROM_DATAPATHS_201;
UNWINDOWED_202 <= FROM_DATAPATHS_202;
UNWINDOWED_203 <= FROM_DATAPATHS_203;
UNWINDOWED_204 <= FROM_DATAPATHS_204;
UNWINDOWED_205 <= FROM_DATAPATHS_205;
UNWINDOWED_206 <= FROM_DATAPATHS_206;
UNWINDOWED_207 <= FROM_DATAPATHS_207;
UNWINDOWED_208 <= FROM_DATAPATHS_208;
UNWINDOWED_209 <= FROM_DATAPATHS_209;
UNWINDOWED_210 <= FROM_DATAPATHS_210;
UNWINDOWED_211 <= FROM_DATAPATHS_211;
UNWINDOWED_212 <= FROM_DATAPATHS_212;
UNWINDOWED_213 <= FROM_DATAPATHS_213;
UNWINDOWED_214 <= FROM_DATAPATHS_214;
UNWINDOWED_215 <= FROM_DATAPATHS_215;
UNWINDOWED_216 <= FROM_DATAPATHS_216;
UNWINDOWED_217 <= FROM_DATAPATHS_217;
UNWINDOWED_218 <= FROM_DATAPATHS_218;
UNWINDOWED_219 <= FROM_DATAPATHS_219;
UNWINDOWED_220 <= FROM_DATAPATHS_220;
UNWINDOWED_221 <= FROM_DATAPATHS_221;
UNWINDOWED_222 <= FROM_DATAPATHS_222;
UNWINDOWED_223 <= FROM_DATAPATHS_223;
UNWINDOWED_224 <= FROM_DATAPATHS_224;
UNWINDOWED_225 <= FROM_DATAPATHS_225;
UNWINDOWED_226 <= FROM_DATAPATHS_226;
UNWINDOWED_227 <= FROM_DATAPATHS_227;
UNWINDOWED_228 <= FROM_DATAPATHS_228;
UNWINDOWED_229 <= FROM_DATAPATHS_229;
UNWINDOWED_230 <= FROM_DATAPATHS_230;
UNWINDOWED_231 <= FROM_DATAPATHS_231;
UNWINDOWED_232 <= FROM_DATAPATHS_232;
UNWINDOWED_233 <= FROM_DATAPATHS_233;
UNWINDOWED_234 <= FROM_DATAPATHS_234;
UNWINDOWED_235 <= FROM_DATAPATHS_235;
UNWINDOWED_236 <= FROM_DATAPATHS_236;
UNWINDOWED_237 <= FROM_DATAPATHS_237;
UNWINDOWED_238 <= FROM_DATAPATHS_238;
UNWINDOWED_239 <= FROM_DATAPATHS_239;
UNWINDOWED_240 <= FROM_DATAPATHS_240;
UNWINDOWED_241 <= FROM_DATAPATHS_241;
UNWINDOWED_242 <= FROM_DATAPATHS_242;
UNWINDOWED_243 <= FROM_DATAPATHS_243;
UNWINDOWED_244 <= FROM_DATAPATHS_244;
UNWINDOWED_245 <= FROM_DATAPATHS_245;
UNWINDOWED_246 <= FROM_DATAPATHS_246;
UNWINDOWED_247 <= FROM_DATAPATHS_247;
UNWINDOWED_248 <= FROM_DATAPATHS_248;
UNWINDOWED_249 <= FROM_DATAPATHS_249;
UNWINDOWED_250 <= FROM_DATAPATHS_250;
UNWINDOWED_251 <= FROM_DATAPATHS_251;
UNWINDOWED_252 <= FROM_DATAPATHS_252;
UNWINDOWED_253 <= FROM_DATAPATHS_253;
UNWINDOWED_254 <= FROM_DATAPATHS_254;
UNWINDOWED_255 <= FROM_DATAPATHS_255;
UNWINDOWED_256 <= FROM_DATAPATHS_256;
UNWINDOWED_257 <= FROM_DATAPATHS_257;
UNWINDOWED_258 <= FROM_DATAPATHS_258;
UNWINDOWED_259 <= FROM_DATAPATHS_259;
UNWINDOWED_260 <= FROM_DATAPATHS_260;
UNWINDOWED_261 <= FROM_DATAPATHS_261;
UNWINDOWED_262 <= FROM_DATAPATHS_262;
UNWINDOWED_263 <= FROM_DATAPATHS_263;
UNWINDOWED_264 <= FROM_DATAPATHS_264;
UNWINDOWED_265 <= FROM_DATAPATHS_265;
UNWINDOWED_266 <= FROM_DATAPATHS_266;
UNWINDOWED_267 <= FROM_DATAPATHS_267;
UNWINDOWED_268 <= FROM_DATAPATHS_268;
UNWINDOWED_269 <= FROM_DATAPATHS_269;
UNWINDOWED_270 <= FROM_DATAPATHS_270;
UNWINDOWED_271 <= FROM_DATAPATHS_271;
UNWINDOWED_272 <= FROM_DATAPATHS_272;
UNWINDOWED_273 <= FROM_DATAPATHS_273;
UNWINDOWED_274 <= FROM_DATAPATHS_274;
UNWINDOWED_275 <= FROM_DATAPATHS_275;
UNWINDOWED_276 <= FROM_DATAPATHS_276;
UNWINDOWED_277 <= FROM_DATAPATHS_277;
UNWINDOWED_278 <= FROM_DATAPATHS_278;
UNWINDOWED_279 <= FROM_DATAPATHS_279;
UNWINDOWED_280 <= FROM_DATAPATHS_280;
UNWINDOWED_281 <= FROM_DATAPATHS_281;
UNWINDOWED_282 <= FROM_DATAPATHS_282;
UNWINDOWED_283 <= FROM_DATAPATHS_283;
UNWINDOWED_284 <= FROM_DATAPATHS_284;
UNWINDOWED_285 <= FROM_DATAPATHS_285;
UNWINDOWED_286 <= FROM_DATAPATHS_286;
UNWINDOWED_287 <= FROM_DATAPATHS_287;
UNWINDOWED_288 <= FROM_DATAPATHS_288;
UNWINDOWED_289 <= FROM_DATAPATHS_289;
UNWINDOWED_290 <= FROM_DATAPATHS_290;
UNWINDOWED_291 <= FROM_DATAPATHS_291;
UNWINDOWED_292 <= FROM_DATAPATHS_292;
UNWINDOWED_293 <= FROM_DATAPATHS_293;
UNWINDOWED_294 <= FROM_DATAPATHS_294;
UNWINDOWED_295 <= FROM_DATAPATHS_295;
UNWINDOWED_296 <= FROM_DATAPATHS_296;
UNWINDOWED_297 <= FROM_DATAPATHS_297;
UNWINDOWED_298 <= FROM_DATAPATHS_298;
UNWINDOWED_299 <= FROM_DATAPATHS_299;
UNWINDOWED_300 <= FROM_DATAPATHS_300;
UNWINDOWED_301 <= FROM_DATAPATHS_301;
UNWINDOWED_302 <= FROM_DATAPATHS_302;
UNWINDOWED_303 <= FROM_DATAPATHS_303;
UNWINDOWED_304 <= FROM_DATAPATHS_304;
UNWINDOWED_305 <= FROM_DATAPATHS_305;
UNWINDOWED_306 <= FROM_DATAPATHS_306;
UNWINDOWED_307 <= FROM_DATAPATHS_307;
UNWINDOWED_308 <= FROM_DATAPATHS_308;
UNWINDOWED_309 <= FROM_DATAPATHS_309;
UNWINDOWED_310 <= FROM_DATAPATHS_310;
UNWINDOWED_311 <= FROM_DATAPATHS_311;
UNWINDOWED_312 <= FROM_DATAPATHS_312;
UNWINDOWED_313 <= FROM_DATAPATHS_313;
UNWINDOWED_314 <= FROM_DATAPATHS_314;
UNWINDOWED_315 <= FROM_DATAPATHS_315;
UNWINDOWED_316 <= FROM_DATAPATHS_316;
UNWINDOWED_317 <= FROM_DATAPATHS_317;
UNWINDOWED_318 <= FROM_DATAPATHS_318;
UNWINDOWED_319 <= FROM_DATAPATHS_319;
UNWINDOWED_320 <= FROM_DATAPATHS_320;
UNWINDOWED_321 <= FROM_DATAPATHS_321;
UNWINDOWED_322 <= FROM_DATAPATHS_322;
UNWINDOWED_323 <= FROM_DATAPATHS_323;
UNWINDOWED_324 <= FROM_DATAPATHS_324;
UNWINDOWED_325 <= FROM_DATAPATHS_325;
UNWINDOWED_326 <= FROM_DATAPATHS_326;
UNWINDOWED_327 <= FROM_DATAPATHS_327;
UNWINDOWED_328 <= FROM_DATAPATHS_328;
UNWINDOWED_329 <= FROM_DATAPATHS_329;
UNWINDOWED_330 <= FROM_DATAPATHS_330;
UNWINDOWED_331 <= FROM_DATAPATHS_331;
UNWINDOWED_332 <= FROM_DATAPATHS_332;
UNWINDOWED_333 <= FROM_DATAPATHS_333;
UNWINDOWED_334 <= FROM_DATAPATHS_334;
UNWINDOWED_335 <= FROM_DATAPATHS_335;
UNWINDOWED_336 <= FROM_DATAPATHS_336;
UNWINDOWED_337 <= FROM_DATAPATHS_337;
UNWINDOWED_338 <= FROM_DATAPATHS_338;
UNWINDOWED_339 <= FROM_DATAPATHS_339;
UNWINDOWED_340 <= FROM_DATAPATHS_340;
UNWINDOWED_341 <= FROM_DATAPATHS_341;
UNWINDOWED_342 <= FROM_DATAPATHS_342;
UNWINDOWED_343 <= FROM_DATAPATHS_343;
UNWINDOWED_344 <= FROM_DATAPATHS_344;
UNWINDOWED_345 <= FROM_DATAPATHS_345;
UNWINDOWED_346 <= FROM_DATAPATHS_346;
UNWINDOWED_347 <= FROM_DATAPATHS_347;
UNWINDOWED_348 <= FROM_DATAPATHS_348;
UNWINDOWED_349 <= FROM_DATAPATHS_349;
UNWINDOWED_350 <= FROM_DATAPATHS_350;
UNWINDOWED_351 <= FROM_DATAPATHS_351;
UNWINDOWED_352 <= FROM_DATAPATHS_352;
UNWINDOWED_353 <= FROM_DATAPATHS_353;
UNWINDOWED_354 <= FROM_DATAPATHS_354;
UNWINDOWED_355 <= FROM_DATAPATHS_355;
UNWINDOWED_356 <= FROM_DATAPATHS_356;
UNWINDOWED_357 <= FROM_DATAPATHS_357;
UNWINDOWED_358 <= FROM_DATAPATHS_358;
UNWINDOWED_359 <= FROM_DATAPATHS_359;
UNWINDOWED_360 <= FROM_DATAPATHS_360;
UNWINDOWED_361 <= FROM_DATAPATHS_361;
UNWINDOWED_362 <= FROM_DATAPATHS_362;
UNWINDOWED_363 <= FROM_DATAPATHS_363;
UNWINDOWED_364 <= FROM_DATAPATHS_364;
UNWINDOWED_365 <= FROM_DATAPATHS_365;
UNWINDOWED_366 <= FROM_DATAPATHS_366;
UNWINDOWED_367 <= FROM_DATAPATHS_367;
UNWINDOWED_368 <= FROM_DATAPATHS_368;
UNWINDOWED_369 <= FROM_DATAPATHS_369;
UNWINDOWED_370 <= FROM_DATAPATHS_370;
UNWINDOWED_371 <= FROM_DATAPATHS_371;
UNWINDOWED_372 <= FROM_DATAPATHS_372;
UNWINDOWED_373 <= FROM_DATAPATHS_373;
UNWINDOWED_374 <= FROM_DATAPATHS_374;
UNWINDOWED_375 <= FROM_DATAPATHS_375;
UNWINDOWED_376 <= FROM_DATAPATHS_376;
UNWINDOWED_377 <= FROM_DATAPATHS_377;
UNWINDOWED_378 <= FROM_DATAPATHS_378;
UNWINDOWED_379 <= FROM_DATAPATHS_379;
UNWINDOWED_380 <= FROM_DATAPATHS_380;
UNWINDOWED_381 <= FROM_DATAPATHS_381;
UNWINDOWED_382 <= FROM_DATAPATHS_382;
UNWINDOWED_383 <= FROM_DATAPATHS_383;
UNWINDOWED_384 <= FROM_DATAPATHS_384;
UNWINDOWED_385 <= FROM_DATAPATHS_385;
UNWINDOWED_386 <= FROM_DATAPATHS_386;
UNWINDOWED_387 <= FROM_DATAPATHS_387;
UNWINDOWED_388 <= FROM_DATAPATHS_388;
UNWINDOWED_389 <= FROM_DATAPATHS_389;
UNWINDOWED_390 <= FROM_DATAPATHS_390;
UNWINDOWED_391 <= FROM_DATAPATHS_391;
UNWINDOWED_392 <= FROM_DATAPATHS_392;
UNWINDOWED_393 <= FROM_DATAPATHS_393;
UNWINDOWED_394 <= FROM_DATAPATHS_394;
UNWINDOWED_395 <= FROM_DATAPATHS_395;
UNWINDOWED_396 <= FROM_DATAPATHS_396;
UNWINDOWED_397 <= FROM_DATAPATHS_397;
UNWINDOWED_398 <= FROM_DATAPATHS_398;
UNWINDOWED_399 <= FROM_DATAPATHS_399;
UNWINDOWED_400 <= FROM_DATAPATHS_400;
UNWINDOWED_401 <= FROM_DATAPATHS_401;
UNWINDOWED_402 <= FROM_DATAPATHS_402;
UNWINDOWED_403 <= FROM_DATAPATHS_403;
UNWINDOWED_404 <= FROM_DATAPATHS_404;
UNWINDOWED_405 <= FROM_DATAPATHS_405;
UNWINDOWED_406 <= FROM_DATAPATHS_406;
UNWINDOWED_407 <= FROM_DATAPATHS_407;
UNWINDOWED_408 <= FROM_DATAPATHS_408;
UNWINDOWED_409 <= FROM_DATAPATHS_409;
UNWINDOWED_410 <= FROM_DATAPATHS_410;
UNWINDOWED_411 <= FROM_DATAPATHS_411;
UNWINDOWED_412 <= FROM_DATAPATHS_412;
UNWINDOWED_413 <= FROM_DATAPATHS_413;
UNWINDOWED_414 <= FROM_DATAPATHS_414;
UNWINDOWED_415 <= FROM_DATAPATHS_415;
UNWINDOWED_416 <= FROM_DATAPATHS_416;
UNWINDOWED_417 <= FROM_DATAPATHS_417;
UNWINDOWED_418 <= FROM_DATAPATHS_418;
UNWINDOWED_419 <= FROM_DATAPATHS_419;
UNWINDOWED_420 <= FROM_DATAPATHS_420;
UNWINDOWED_421 <= FROM_DATAPATHS_421;
UNWINDOWED_422 <= FROM_DATAPATHS_422;
UNWINDOWED_423 <= FROM_DATAPATHS_423;
UNWINDOWED_424 <= FROM_DATAPATHS_424;
UNWINDOWED_425 <= FROM_DATAPATHS_425;
UNWINDOWED_426 <= FROM_DATAPATHS_426;
UNWINDOWED_427 <= FROM_DATAPATHS_427;
UNWINDOWED_428 <= FROM_DATAPATHS_428;
UNWINDOWED_429 <= FROM_DATAPATHS_429;
UNWINDOWED_430 <= FROM_DATAPATHS_430;
UNWINDOWED_431 <= FROM_DATAPATHS_431;
UNWINDOWED_432 <= FROM_DATAPATHS_432;
UNWINDOWED_433 <= FROM_DATAPATHS_433;
UNWINDOWED_434 <= FROM_DATAPATHS_434;
UNWINDOWED_435 <= FROM_DATAPATHS_435;
UNWINDOWED_436 <= FROM_DATAPATHS_436;
UNWINDOWED_437 <= FROM_DATAPATHS_437;
UNWINDOWED_438 <= FROM_DATAPATHS_438;
UNWINDOWED_439 <= FROM_DATAPATHS_439;
UNWINDOWED_440 <= FROM_DATAPATHS_440;
UNWINDOWED_441 <= FROM_DATAPATHS_441;
UNWINDOWED_442 <= FROM_DATAPATHS_442;
UNWINDOWED_443 <= FROM_DATAPATHS_443;
UNWINDOWED_444 <= FROM_DATAPATHS_444;
UNWINDOWED_445 <= FROM_DATAPATHS_445;
UNWINDOWED_446 <= FROM_DATAPATHS_446;
UNWINDOWED_447 <= FROM_DATAPATHS_447;
UNWINDOWED_448 <= FROM_DATAPATHS_448;
UNWINDOWED_449 <= FROM_DATAPATHS_449;
UNWINDOWED_450 <= FROM_DATAPATHS_450;
UNWINDOWED_451 <= FROM_DATAPATHS_451;
UNWINDOWED_452 <= FROM_DATAPATHS_452;
UNWINDOWED_453 <= FROM_DATAPATHS_453;
UNWINDOWED_454 <= FROM_DATAPATHS_454;
UNWINDOWED_455 <= FROM_DATAPATHS_455;
UNWINDOWED_456 <= FROM_DATAPATHS_456;
UNWINDOWED_457 <= FROM_DATAPATHS_457;
UNWINDOWED_458 <= FROM_DATAPATHS_458;
UNWINDOWED_459 <= FROM_DATAPATHS_459;
UNWINDOWED_460 <= FROM_DATAPATHS_460;
UNWINDOWED_461 <= FROM_DATAPATHS_461;
UNWINDOWED_462 <= FROM_DATAPATHS_462;
UNWINDOWED_463 <= FROM_DATAPATHS_463;
UNWINDOWED_464 <= FROM_DATAPATHS_464;
UNWINDOWED_465 <= FROM_DATAPATHS_465;
UNWINDOWED_466 <= FROM_DATAPATHS_466;
UNWINDOWED_467 <= FROM_DATAPATHS_467;
UNWINDOWED_468 <= FROM_DATAPATHS_468;
UNWINDOWED_469 <= FROM_DATAPATHS_469;
UNWINDOWED_470 <= FROM_DATAPATHS_470;
UNWINDOWED_471 <= FROM_DATAPATHS_471;
UNWINDOWED_472 <= FROM_DATAPATHS_472;
UNWINDOWED_473 <= FROM_DATAPATHS_473;
UNWINDOWED_474 <= FROM_DATAPATHS_474;
UNWINDOWED_475 <= FROM_DATAPATHS_475;
UNWINDOWED_476 <= FROM_DATAPATHS_476;
UNWINDOWED_477 <= FROM_DATAPATHS_477;
UNWINDOWED_478 <= FROM_DATAPATHS_478;
UNWINDOWED_479 <= FROM_DATAPATHS_479;
UNWINDOWED_480 <= FROM_DATAPATHS_480;
UNWINDOWED_481 <= FROM_DATAPATHS_481;
UNWINDOWED_482 <= FROM_DATAPATHS_482;
UNWINDOWED_483 <= FROM_DATAPATHS_483;
UNWINDOWED_484 <= FROM_DATAPATHS_484;
UNWINDOWED_485 <= FROM_DATAPATHS_485;
UNWINDOWED_486 <= FROM_DATAPATHS_486;
UNWINDOWED_487 <= FROM_DATAPATHS_487;
UNWINDOWED_488 <= FROM_DATAPATHS_488;
UNWINDOWED_489 <= FROM_DATAPATHS_489;
UNWINDOWED_490 <= FROM_DATAPATHS_490;
UNWINDOWED_491 <= FROM_DATAPATHS_491;
UNWINDOWED_492 <= FROM_DATAPATHS_492;
UNWINDOWED_493 <= FROM_DATAPATHS_493;
UNWINDOWED_494 <= FROM_DATAPATHS_494;
UNWINDOWED_495 <= FROM_DATAPATHS_495;
UNWINDOWED_496 <= FROM_DATAPATHS_496;
UNWINDOWED_497 <= FROM_DATAPATHS_497;
UNWINDOWED_498 <= FROM_DATAPATHS_498;
UNWINDOWED_499 <= FROM_DATAPATHS_499;
UNWINDOWED_500 <= FROM_DATAPATHS_500;
UNWINDOWED_501 <= FROM_DATAPATHS_501;
UNWINDOWED_502 <= FROM_DATAPATHS_502;
UNWINDOWED_503 <= FROM_DATAPATHS_503;
UNWINDOWED_504 <= FROM_DATAPATHS_504;
UNWINDOWED_505 <= FROM_DATAPATHS_505;
UNWINDOWED_506 <= FROM_DATAPATHS_506;
UNWINDOWED_507 <= FROM_DATAPATHS_507;
UNWINDOWED_508 <= FROM_DATAPATHS_508;
UNWINDOWED_509 <= FROM_DATAPATHS_509;
UNWINDOWED_510 <= FROM_DATAPATHS_510;
UNWINDOWED_511 <= FROM_DATAPATHS_511;
UNWINDOWED_512 <= FROM_DATAPATHS_512;
UNWINDOWED_513 <= FROM_DATAPATHS_513;
UNWINDOWED_514 <= FROM_DATAPATHS_514;
UNWINDOWED_515 <= FROM_DATAPATHS_515;
UNWINDOWED_516 <= FROM_DATAPATHS_516;
UNWINDOWED_517 <= FROM_DATAPATHS_517;
UNWINDOWED_518 <= FROM_DATAPATHS_518;
UNWINDOWED_519 <= FROM_DATAPATHS_519;
UNWINDOWED_520 <= FROM_DATAPATHS_520;
UNWINDOWED_521 <= FROM_DATAPATHS_521;
UNWINDOWED_522 <= FROM_DATAPATHS_522;
UNWINDOWED_523 <= FROM_DATAPATHS_523;
UNWINDOWED_524 <= FROM_DATAPATHS_524;
UNWINDOWED_525 <= FROM_DATAPATHS_525;
UNWINDOWED_526 <= FROM_DATAPATHS_526;
UNWINDOWED_527 <= FROM_DATAPATHS_527;
UNWINDOWED_528 <= FROM_DATAPATHS_528;
UNWINDOWED_529 <= FROM_DATAPATHS_529;
UNWINDOWED_530 <= FROM_DATAPATHS_530;
UNWINDOWED_531 <= FROM_DATAPATHS_531;
UNWINDOWED_532 <= FROM_DATAPATHS_532;
UNWINDOWED_533 <= FROM_DATAPATHS_533;
UNWINDOWED_534 <= FROM_DATAPATHS_534;
UNWINDOWED_535 <= FROM_DATAPATHS_535;
UNWINDOWED_536 <= FROM_DATAPATHS_536;
UNWINDOWED_537 <= FROM_DATAPATHS_537;
UNWINDOWED_538 <= FROM_DATAPATHS_538;
UNWINDOWED_539 <= FROM_DATAPATHS_539;
UNWINDOWED_540 <= FROM_DATAPATHS_540;
UNWINDOWED_541 <= FROM_DATAPATHS_541;
UNWINDOWED_542 <= FROM_DATAPATHS_542;
UNWINDOWED_543 <= FROM_DATAPATHS_543;
UNWINDOWED_544 <= FROM_DATAPATHS_544;
UNWINDOWED_545 <= FROM_DATAPATHS_545;
UNWINDOWED_546 <= FROM_DATAPATHS_546;
UNWINDOWED_547 <= FROM_DATAPATHS_547;
UNWINDOWED_548 <= FROM_DATAPATHS_548;
UNWINDOWED_549 <= FROM_DATAPATHS_549;
UNWINDOWED_550 <= FROM_DATAPATHS_550;
UNWINDOWED_551 <= FROM_DATAPATHS_551;
UNWINDOWED_552 <= FROM_DATAPATHS_552;
UNWINDOWED_553 <= FROM_DATAPATHS_553;
UNWINDOWED_554 <= FROM_DATAPATHS_554;
UNWINDOWED_555 <= FROM_DATAPATHS_555;
UNWINDOWED_556 <= FROM_DATAPATHS_556;
UNWINDOWED_557 <= FROM_DATAPATHS_557;
UNWINDOWED_558 <= FROM_DATAPATHS_558;
UNWINDOWED_559 <= FROM_DATAPATHS_559;
UNWINDOWED_560 <= FROM_DATAPATHS_560;
UNWINDOWED_561 <= FROM_DATAPATHS_561;
UNWINDOWED_562 <= FROM_DATAPATHS_562;
UNWINDOWED_563 <= FROM_DATAPATHS_563;
UNWINDOWED_564 <= FROM_DATAPATHS_564;
UNWINDOWED_565 <= FROM_DATAPATHS_565;
UNWINDOWED_566 <= FROM_DATAPATHS_566;
UNWINDOWED_567 <= FROM_DATAPATHS_567;
UNWINDOWED_568 <= FROM_DATAPATHS_568;
UNWINDOWED_569 <= FROM_DATAPATHS_569;
UNWINDOWED_570 <= FROM_DATAPATHS_570;
UNWINDOWED_571 <= FROM_DATAPATHS_571;
UNWINDOWED_572 <= FROM_DATAPATHS_572;
UNWINDOWED_573 <= FROM_DATAPATHS_573;
UNWINDOWED_574 <= FROM_DATAPATHS_574;
UNWINDOWED_575 <= FROM_DATAPATHS_575;
UNWINDOWED_576 <= FROM_DATAPATHS_576;
UNWINDOWED_577 <= FROM_DATAPATHS_577;
UNWINDOWED_578 <= FROM_DATAPATHS_578;
UNWINDOWED_579 <= FROM_DATAPATHS_579;
UNWINDOWED_580 <= FROM_DATAPATHS_580;
UNWINDOWED_581 <= FROM_DATAPATHS_581;
UNWINDOWED_582 <= FROM_DATAPATHS_582;
UNWINDOWED_583 <= FROM_DATAPATHS_583;
UNWINDOWED_584 <= FROM_DATAPATHS_584;
UNWINDOWED_585 <= FROM_DATAPATHS_585;
UNWINDOWED_586 <= FROM_DATAPATHS_586;
UNWINDOWED_587 <= FROM_DATAPATHS_587;
UNWINDOWED_588 <= FROM_DATAPATHS_588;
UNWINDOWED_589 <= FROM_DATAPATHS_589;
UNWINDOWED_590 <= FROM_DATAPATHS_590;
UNWINDOWED_591 <= FROM_DATAPATHS_591;
UNWINDOWED_592 <= FROM_DATAPATHS_592;
UNWINDOWED_593 <= FROM_DATAPATHS_593;
UNWINDOWED_594 <= FROM_DATAPATHS_594;
UNWINDOWED_595 <= FROM_DATAPATHS_595;
UNWINDOWED_596 <= FROM_DATAPATHS_596;
UNWINDOWED_597 <= FROM_DATAPATHS_597;
UNWINDOWED_598 <= FROM_DATAPATHS_598;
UNWINDOWED_599 <= FROM_DATAPATHS_599;
UNWINDOWED_600 <= FROM_DATAPATHS_600;
UNWINDOWED_601 <= FROM_DATAPATHS_601;
UNWINDOWED_602 <= FROM_DATAPATHS_602;
UNWINDOWED_603 <= FROM_DATAPATHS_603;
UNWINDOWED_604 <= FROM_DATAPATHS_604;
UNWINDOWED_605 <= FROM_DATAPATHS_605;
UNWINDOWED_606 <= FROM_DATAPATHS_606;
UNWINDOWED_607 <= FROM_DATAPATHS_607;
UNWINDOWED_608 <= FROM_DATAPATHS_608;
UNWINDOWED_609 <= FROM_DATAPATHS_609;
UNWINDOWED_610 <= FROM_DATAPATHS_610;
UNWINDOWED_611 <= FROM_DATAPATHS_611;
UNWINDOWED_612 <= FROM_DATAPATHS_612;
UNWINDOWED_613 <= FROM_DATAPATHS_613;
UNWINDOWED_614 <= FROM_DATAPATHS_614;
UNWINDOWED_615 <= FROM_DATAPATHS_615;
UNWINDOWED_616 <= FROM_DATAPATHS_616;
UNWINDOWED_617 <= FROM_DATAPATHS_617;
UNWINDOWED_618 <= FROM_DATAPATHS_618;
UNWINDOWED_619 <= FROM_DATAPATHS_619;
UNWINDOWED_620 <= FROM_DATAPATHS_620;
UNWINDOWED_621 <= FROM_DATAPATHS_621;
UNWINDOWED_622 <= FROM_DATAPATHS_622;
UNWINDOWED_623 <= FROM_DATAPATHS_623;
UNWINDOWED_624 <= FROM_DATAPATHS_624;
UNWINDOWED_625 <= FROM_DATAPATHS_625;
UNWINDOWED_626 <= FROM_DATAPATHS_626;
UNWINDOWED_627 <= FROM_DATAPATHS_627;
UNWINDOWED_628 <= FROM_DATAPATHS_628;
UNWINDOWED_629 <= FROM_DATAPATHS_629;
UNWINDOWED_630 <= FROM_DATAPATHS_630;
UNWINDOWED_631 <= FROM_DATAPATHS_631;
UNWINDOWED_632 <= FROM_DATAPATHS_632;
UNWINDOWED_633 <= FROM_DATAPATHS_633;
UNWINDOWED_634 <= FROM_DATAPATHS_634;
UNWINDOWED_635 <= FROM_DATAPATHS_635;
UNWINDOWED_636 <= FROM_DATAPATHS_636;
UNWINDOWED_637 <= FROM_DATAPATHS_637;
UNWINDOWED_638 <= FROM_DATAPATHS_638;
UNWINDOWED_639 <= FROM_DATAPATHS_639;
UNWINDOWED_640 <= FROM_DATAPATHS_640;
UNWINDOWED_641 <= FROM_DATAPATHS_641;
UNWINDOWED_642 <= FROM_DATAPATHS_642;
UNWINDOWED_643 <= FROM_DATAPATHS_643;
UNWINDOWED_644 <= FROM_DATAPATHS_644;
UNWINDOWED_645 <= FROM_DATAPATHS_645;
UNWINDOWED_646 <= FROM_DATAPATHS_646;
UNWINDOWED_647 <= FROM_DATAPATHS_647;
UNWINDOWED_648 <= FROM_DATAPATHS_648;
UNWINDOWED_649 <= FROM_DATAPATHS_649;
UNWINDOWED_650 <= FROM_DATAPATHS_650;
UNWINDOWED_651 <= FROM_DATAPATHS_651;
UNWINDOWED_652 <= FROM_DATAPATHS_652;
UNWINDOWED_653 <= FROM_DATAPATHS_653;
UNWINDOWED_654 <= FROM_DATAPATHS_654;
UNWINDOWED_655 <= FROM_DATAPATHS_655;
UNWINDOWED_656 <= FROM_DATAPATHS_656;
UNWINDOWED_657 <= FROM_DATAPATHS_657;
UNWINDOWED_658 <= FROM_DATAPATHS_658;
UNWINDOWED_659 <= FROM_DATAPATHS_659;
UNWINDOWED_660 <= FROM_DATAPATHS_660;
UNWINDOWED_661 <= FROM_DATAPATHS_661;
UNWINDOWED_662 <= FROM_DATAPATHS_662;
UNWINDOWED_663 <= FROM_DATAPATHS_663;
UNWINDOWED_664 <= FROM_DATAPATHS_664;
UNWINDOWED_665 <= FROM_DATAPATHS_665;
UNWINDOWED_666 <= FROM_DATAPATHS_666;
UNWINDOWED_667 <= FROM_DATAPATHS_667;
UNWINDOWED_668 <= FROM_DATAPATHS_668;
UNWINDOWED_669 <= FROM_DATAPATHS_669;
UNWINDOWED_670 <= FROM_DATAPATHS_670;
UNWINDOWED_671 <= FROM_DATAPATHS_671;
UNWINDOWED_672 <= FROM_DATAPATHS_672;
UNWINDOWED_673 <= FROM_DATAPATHS_673;
UNWINDOWED_674 <= FROM_DATAPATHS_674;
UNWINDOWED_675 <= FROM_DATAPATHS_675;
UNWINDOWED_676 <= FROM_DATAPATHS_676;
UNWINDOWED_677 <= FROM_DATAPATHS_677;
UNWINDOWED_678 <= FROM_DATAPATHS_678;
UNWINDOWED_679 <= FROM_DATAPATHS_679;
UNWINDOWED_680 <= FROM_DATAPATHS_680;
UNWINDOWED_681 <= FROM_DATAPATHS_681;
UNWINDOWED_682 <= FROM_DATAPATHS_682;
UNWINDOWED_683 <= FROM_DATAPATHS_683;
UNWINDOWED_684 <= FROM_DATAPATHS_684;
UNWINDOWED_685 <= FROM_DATAPATHS_685;
UNWINDOWED_686 <= FROM_DATAPATHS_686;
UNWINDOWED_687 <= FROM_DATAPATHS_687;
UNWINDOWED_688 <= FROM_DATAPATHS_688;
UNWINDOWED_689 <= FROM_DATAPATHS_689;
UNWINDOWED_690 <= FROM_DATAPATHS_690;
UNWINDOWED_691 <= FROM_DATAPATHS_691;
UNWINDOWED_692 <= FROM_DATAPATHS_692;
UNWINDOWED_693 <= FROM_DATAPATHS_693;
UNWINDOWED_694 <= FROM_DATAPATHS_694;
UNWINDOWED_695 <= FROM_DATAPATHS_695;
UNWINDOWED_696 <= FROM_DATAPATHS_696;
UNWINDOWED_697 <= FROM_DATAPATHS_697;
UNWINDOWED_698 <= FROM_DATAPATHS_698;
UNWINDOWED_699 <= FROM_DATAPATHS_699;
UNWINDOWED_700 <= FROM_DATAPATHS_700;
UNWINDOWED_701 <= FROM_DATAPATHS_701;
UNWINDOWED_702 <= FROM_DATAPATHS_702;
UNWINDOWED_703 <= FROM_DATAPATHS_703;
UNWINDOWED_704 <= FROM_DATAPATHS_704;
UNWINDOWED_705 <= FROM_DATAPATHS_705;
UNWINDOWED_706 <= FROM_DATAPATHS_706;
UNWINDOWED_707 <= FROM_DATAPATHS_707;
UNWINDOWED_708 <= FROM_DATAPATHS_708;
UNWINDOWED_709 <= FROM_DATAPATHS_709;
UNWINDOWED_710 <= FROM_DATAPATHS_710;
UNWINDOWED_711 <= FROM_DATAPATHS_711;
UNWINDOWED_712 <= FROM_DATAPATHS_712;
UNWINDOWED_713 <= FROM_DATAPATHS_713;
UNWINDOWED_714 <= FROM_DATAPATHS_714;
UNWINDOWED_715 <= FROM_DATAPATHS_715;
UNWINDOWED_716 <= FROM_DATAPATHS_716;
UNWINDOWED_717 <= FROM_DATAPATHS_717;
UNWINDOWED_718 <= FROM_DATAPATHS_718;
UNWINDOWED_719 <= FROM_DATAPATHS_719;
UNWINDOWED_720 <= FROM_DATAPATHS_720;
UNWINDOWED_721 <= FROM_DATAPATHS_721;
UNWINDOWED_722 <= FROM_DATAPATHS_722;
UNWINDOWED_723 <= FROM_DATAPATHS_723;
UNWINDOWED_724 <= FROM_DATAPATHS_724;
UNWINDOWED_725 <= FROM_DATAPATHS_725;
UNWINDOWED_726 <= FROM_DATAPATHS_726;
UNWINDOWED_727 <= FROM_DATAPATHS_727;
UNWINDOWED_728 <= FROM_DATAPATHS_728;
UNWINDOWED_729 <= FROM_DATAPATHS_729;
UNWINDOWED_730 <= FROM_DATAPATHS_730;
UNWINDOWED_731 <= FROM_DATAPATHS_731;
UNWINDOWED_732 <= FROM_DATAPATHS_732;
UNWINDOWED_733 <= FROM_DATAPATHS_733;
UNWINDOWED_734 <= FROM_DATAPATHS_734;
UNWINDOWED_735 <= FROM_DATAPATHS_735;
UNWINDOWED_736 <= FROM_DATAPATHS_736;
UNWINDOWED_737 <= FROM_DATAPATHS_737;
UNWINDOWED_738 <= FROM_DATAPATHS_738;
UNWINDOWED_739 <= FROM_DATAPATHS_739;
UNWINDOWED_740 <= FROM_DATAPATHS_740;
UNWINDOWED_741 <= FROM_DATAPATHS_741;
UNWINDOWED_742 <= FROM_DATAPATHS_742;
UNWINDOWED_743 <= FROM_DATAPATHS_743;
UNWINDOWED_744 <= FROM_DATAPATHS_744;
UNWINDOWED_745 <= FROM_DATAPATHS_745;
UNWINDOWED_746 <= FROM_DATAPATHS_746;
UNWINDOWED_747 <= FROM_DATAPATHS_747;
UNWINDOWED_748 <= FROM_DATAPATHS_748;
UNWINDOWED_749 <= FROM_DATAPATHS_749;
UNWINDOWED_750 <= FROM_DATAPATHS_750;
UNWINDOWED_751 <= FROM_DATAPATHS_751;
UNWINDOWED_752 <= FROM_DATAPATHS_752;
UNWINDOWED_753 <= FROM_DATAPATHS_753;
UNWINDOWED_754 <= FROM_DATAPATHS_754;
UNWINDOWED_755 <= FROM_DATAPATHS_755;
UNWINDOWED_756 <= FROM_DATAPATHS_756;
UNWINDOWED_757 <= FROM_DATAPATHS_757;
UNWINDOWED_758 <= FROM_DATAPATHS_758;
UNWINDOWED_759 <= FROM_DATAPATHS_759;
UNWINDOWED_760 <= FROM_DATAPATHS_760;
UNWINDOWED_761 <= FROM_DATAPATHS_761;
UNWINDOWED_762 <= FROM_DATAPATHS_762;
UNWINDOWED_763 <= FROM_DATAPATHS_763;
UNWINDOWED_764 <= FROM_DATAPATHS_764;
UNWINDOWED_765 <= FROM_DATAPATHS_765;
UNWINDOWED_766 <= FROM_DATAPATHS_766;
UNWINDOWED_767 <= FROM_DATAPATHS_767;
UNWINDOWED_768 <= FROM_DATAPATHS_768;
UNWINDOWED_769 <= FROM_DATAPATHS_769;
UNWINDOWED_770 <= FROM_DATAPATHS_770;
UNWINDOWED_771 <= FROM_DATAPATHS_771;
UNWINDOWED_772 <= FROM_DATAPATHS_772;
UNWINDOWED_773 <= FROM_DATAPATHS_773;
UNWINDOWED_774 <= FROM_DATAPATHS_774;
UNWINDOWED_775 <= FROM_DATAPATHS_775;
UNWINDOWED_776 <= FROM_DATAPATHS_776;
UNWINDOWED_777 <= FROM_DATAPATHS_777;
UNWINDOWED_778 <= FROM_DATAPATHS_778;
UNWINDOWED_779 <= FROM_DATAPATHS_779;
UNWINDOWED_780 <= FROM_DATAPATHS_780;
UNWINDOWED_781 <= FROM_DATAPATHS_781;
UNWINDOWED_782 <= FROM_DATAPATHS_782;
UNWINDOWED_783 <= FROM_DATAPATHS_783;
UNWINDOWED_784 <= FROM_DATAPATHS_784;
UNWINDOWED_785 <= FROM_DATAPATHS_785;
UNWINDOWED_786 <= FROM_DATAPATHS_786;
UNWINDOWED_787 <= FROM_DATAPATHS_787;
UNWINDOWED_788 <= FROM_DATAPATHS_788;
UNWINDOWED_789 <= FROM_DATAPATHS_789;
UNWINDOWED_790 <= FROM_DATAPATHS_790;
UNWINDOWED_791 <= FROM_DATAPATHS_791;
UNWINDOWED_792 <= FROM_DATAPATHS_792;
UNWINDOWED_793 <= FROM_DATAPATHS_793;
UNWINDOWED_794 <= FROM_DATAPATHS_794;
UNWINDOWED_795 <= FROM_DATAPATHS_795;
UNWINDOWED_796 <= FROM_DATAPATHS_796;
UNWINDOWED_797 <= FROM_DATAPATHS_797;
UNWINDOWED_798 <= FROM_DATAPATHS_798;
UNWINDOWED_799 <= FROM_DATAPATHS_799;
UNWINDOWED_800 <= FROM_DATAPATHS_800;
UNWINDOWED_801 <= FROM_DATAPATHS_801;
UNWINDOWED_802 <= FROM_DATAPATHS_802;
UNWINDOWED_803 <= FROM_DATAPATHS_803;
UNWINDOWED_804 <= FROM_DATAPATHS_804;
UNWINDOWED_805 <= FROM_DATAPATHS_805;
UNWINDOWED_806 <= FROM_DATAPATHS_806;
UNWINDOWED_807 <= FROM_DATAPATHS_807;
UNWINDOWED_808 <= FROM_DATAPATHS_808;
UNWINDOWED_809 <= FROM_DATAPATHS_809;
UNWINDOWED_810 <= FROM_DATAPATHS_810;
UNWINDOWED_811 <= FROM_DATAPATHS_811;
UNWINDOWED_812 <= FROM_DATAPATHS_812;
UNWINDOWED_813 <= FROM_DATAPATHS_813;
UNWINDOWED_814 <= FROM_DATAPATHS_814;
UNWINDOWED_815 <= FROM_DATAPATHS_815;
UNWINDOWED_816 <= FROM_DATAPATHS_816;
UNWINDOWED_817 <= FROM_DATAPATHS_817;
UNWINDOWED_818 <= FROM_DATAPATHS_818;
UNWINDOWED_819 <= FROM_DATAPATHS_819;
UNWINDOWED_820 <= FROM_DATAPATHS_820;
UNWINDOWED_821 <= FROM_DATAPATHS_821;
UNWINDOWED_822 <= FROM_DATAPATHS_822;
UNWINDOWED_823 <= FROM_DATAPATHS_823;
UNWINDOWED_824 <= FROM_DATAPATHS_824;
UNWINDOWED_825 <= FROM_DATAPATHS_825;
UNWINDOWED_826 <= FROM_DATAPATHS_826;
UNWINDOWED_827 <= FROM_DATAPATHS_827;
UNWINDOWED_828 <= FROM_DATAPATHS_828;
UNWINDOWED_829 <= FROM_DATAPATHS_829;
UNWINDOWED_830 <= FROM_DATAPATHS_830;
UNWINDOWED_831 <= FROM_DATAPATHS_831;
UNWINDOWED_832 <= FROM_DATAPATHS_832;
UNWINDOWED_833 <= FROM_DATAPATHS_833;
UNWINDOWED_834 <= FROM_DATAPATHS_834;
UNWINDOWED_835 <= FROM_DATAPATHS_835;
UNWINDOWED_836 <= FROM_DATAPATHS_836;
UNWINDOWED_837 <= FROM_DATAPATHS_837;
UNWINDOWED_838 <= FROM_DATAPATHS_838;
UNWINDOWED_839 <= FROM_DATAPATHS_839;
UNWINDOWED_840 <= FROM_DATAPATHS_840;
UNWINDOWED_841 <= FROM_DATAPATHS_841;
UNWINDOWED_842 <= FROM_DATAPATHS_842;
UNWINDOWED_843 <= FROM_DATAPATHS_843;
UNWINDOWED_844 <= FROM_DATAPATHS_844;
UNWINDOWED_845 <= FROM_DATAPATHS_845;
UNWINDOWED_846 <= FROM_DATAPATHS_846;
UNWINDOWED_847 <= FROM_DATAPATHS_847;
UNWINDOWED_848 <= FROM_DATAPATHS_848;
UNWINDOWED_849 <= FROM_DATAPATHS_849;
UNWINDOWED_850 <= FROM_DATAPATHS_850;
UNWINDOWED_851 <= FROM_DATAPATHS_851;
UNWINDOWED_852 <= FROM_DATAPATHS_852;
UNWINDOWED_853 <= FROM_DATAPATHS_853;
UNWINDOWED_854 <= FROM_DATAPATHS_854;
UNWINDOWED_855 <= FROM_DATAPATHS_855;
UNWINDOWED_856 <= FROM_DATAPATHS_856;
UNWINDOWED_857 <= FROM_DATAPATHS_857;
UNWINDOWED_858 <= FROM_DATAPATHS_858;
UNWINDOWED_859 <= FROM_DATAPATHS_859;
UNWINDOWED_860 <= FROM_DATAPATHS_860;
UNWINDOWED_861 <= FROM_DATAPATHS_861;
UNWINDOWED_862 <= FROM_DATAPATHS_862;
UNWINDOWED_863 <= FROM_DATAPATHS_863;
UNWINDOWED_864 <= FROM_DATAPATHS_864;
UNWINDOWED_865 <= FROM_DATAPATHS_865;
UNWINDOWED_866 <= FROM_DATAPATHS_866;
UNWINDOWED_867 <= FROM_DATAPATHS_867;
UNWINDOWED_868 <= FROM_DATAPATHS_868;
UNWINDOWED_869 <= FROM_DATAPATHS_869;
UNWINDOWED_870 <= FROM_DATAPATHS_870;
UNWINDOWED_871 <= FROM_DATAPATHS_871;
UNWINDOWED_872 <= FROM_DATAPATHS_872;
UNWINDOWED_873 <= FROM_DATAPATHS_873;
UNWINDOWED_874 <= FROM_DATAPATHS_874;
UNWINDOWED_875 <= FROM_DATAPATHS_875;
UNWINDOWED_876 <= FROM_DATAPATHS_876;
UNWINDOWED_877 <= FROM_DATAPATHS_877;
UNWINDOWED_878 <= FROM_DATAPATHS_878;
UNWINDOWED_879 <= FROM_DATAPATHS_879;
UNWINDOWED_880 <= FROM_DATAPATHS_880;
UNWINDOWED_881 <= FROM_DATAPATHS_881;
UNWINDOWED_882 <= FROM_DATAPATHS_882;
UNWINDOWED_883 <= FROM_DATAPATHS_883;
UNWINDOWED_884 <= FROM_DATAPATHS_884;
UNWINDOWED_885 <= FROM_DATAPATHS_885;
UNWINDOWED_886 <= FROM_DATAPATHS_886;
UNWINDOWED_887 <= FROM_DATAPATHS_887;
UNWINDOWED_888 <= FROM_DATAPATHS_888;
UNWINDOWED_889 <= FROM_DATAPATHS_889;
UNWINDOWED_890 <= FROM_DATAPATHS_890;
UNWINDOWED_891 <= FROM_DATAPATHS_891;
UNWINDOWED_892 <= FROM_DATAPATHS_892;
UNWINDOWED_893 <= FROM_DATAPATHS_893;
UNWINDOWED_894 <= FROM_DATAPATHS_894;
UNWINDOWED_895 <= FROM_DATAPATHS_895;
UNWINDOWED_896 <= FROM_DATAPATHS_896;
UNWINDOWED_897 <= FROM_DATAPATHS_897;
UNWINDOWED_898 <= FROM_DATAPATHS_898;
UNWINDOWED_899 <= FROM_DATAPATHS_899;
UNWINDOWED_900 <= FROM_DATAPATHS_900;
UNWINDOWED_901 <= FROM_DATAPATHS_901;
UNWINDOWED_902 <= FROM_DATAPATHS_902;
UNWINDOWED_903 <= FROM_DATAPATHS_903;
UNWINDOWED_904 <= FROM_DATAPATHS_904;
UNWINDOWED_905 <= FROM_DATAPATHS_905;
UNWINDOWED_906 <= FROM_DATAPATHS_906;
UNWINDOWED_907 <= FROM_DATAPATHS_907;
UNWINDOWED_908 <= FROM_DATAPATHS_908;
UNWINDOWED_909 <= FROM_DATAPATHS_909;
UNWINDOWED_910 <= FROM_DATAPATHS_910;
UNWINDOWED_911 <= FROM_DATAPATHS_911;
UNWINDOWED_912 <= FROM_DATAPATHS_912;
UNWINDOWED_913 <= FROM_DATAPATHS_913;
UNWINDOWED_914 <= FROM_DATAPATHS_914;
UNWINDOWED_915 <= FROM_DATAPATHS_915;
UNWINDOWED_916 <= FROM_DATAPATHS_916;
UNWINDOWED_917 <= FROM_DATAPATHS_917;
UNWINDOWED_918 <= FROM_DATAPATHS_918;
UNWINDOWED_919 <= FROM_DATAPATHS_919;
UNWINDOWED_920 <= FROM_DATAPATHS_920;
UNWINDOWED_921 <= FROM_DATAPATHS_921;
UNWINDOWED_922 <= FROM_DATAPATHS_922;
UNWINDOWED_923 <= FROM_DATAPATHS_923;
UNWINDOWED_924 <= FROM_DATAPATHS_924;
UNWINDOWED_925 <= FROM_DATAPATHS_925;
UNWINDOWED_926 <= FROM_DATAPATHS_926;
UNWINDOWED_927 <= FROM_DATAPATHS_927;
UNWINDOWED_928 <= FROM_DATAPATHS_928;
UNWINDOWED_929 <= FROM_DATAPATHS_929;
UNWINDOWED_930 <= FROM_DATAPATHS_930;
UNWINDOWED_931 <= FROM_DATAPATHS_931;
UNWINDOWED_932 <= FROM_DATAPATHS_932;
UNWINDOWED_933 <= FROM_DATAPATHS_933;
UNWINDOWED_934 <= FROM_DATAPATHS_934;
UNWINDOWED_935 <= FROM_DATAPATHS_935;
UNWINDOWED_936 <= FROM_DATAPATHS_936;
UNWINDOWED_937 <= FROM_DATAPATHS_937;
UNWINDOWED_938 <= FROM_DATAPATHS_938;
UNWINDOWED_939 <= FROM_DATAPATHS_939;
UNWINDOWED_940 <= FROM_DATAPATHS_940;
UNWINDOWED_941 <= FROM_DATAPATHS_941;
UNWINDOWED_942 <= FROM_DATAPATHS_942;
UNWINDOWED_943 <= FROM_DATAPATHS_943;
UNWINDOWED_944 <= FROM_DATAPATHS_944;
UNWINDOWED_945 <= FROM_DATAPATHS_945;
UNWINDOWED_946 <= FROM_DATAPATHS_946;
UNWINDOWED_947 <= FROM_DATAPATHS_947;
UNWINDOWED_948 <= FROM_DATAPATHS_948;
UNWINDOWED_949 <= FROM_DATAPATHS_949;
UNWINDOWED_950 <= FROM_DATAPATHS_950;
UNWINDOWED_951 <= FROM_DATAPATHS_951;
UNWINDOWED_952 <= FROM_DATAPATHS_952;
UNWINDOWED_953 <= FROM_DATAPATHS_953;
UNWINDOWED_954 <= FROM_DATAPATHS_954;
UNWINDOWED_955 <= FROM_DATAPATHS_955;
UNWINDOWED_956 <= FROM_DATAPATHS_956;
UNWINDOWED_957 <= FROM_DATAPATHS_957;
UNWINDOWED_958 <= FROM_DATAPATHS_958;
UNWINDOWED_959 <= FROM_DATAPATHS_959;
UNWINDOWED_960 <= FROM_DATAPATHS_960;
UNWINDOWED_961 <= FROM_DATAPATHS_961;
UNWINDOWED_962 <= FROM_DATAPATHS_962;
UNWINDOWED_963 <= FROM_DATAPATHS_963;
UNWINDOWED_964 <= FROM_DATAPATHS_964;
UNWINDOWED_965 <= FROM_DATAPATHS_965;
UNWINDOWED_966 <= FROM_DATAPATHS_966;
UNWINDOWED_967 <= FROM_DATAPATHS_967;
UNWINDOWED_968 <= FROM_DATAPATHS_968;
UNWINDOWED_969 <= FROM_DATAPATHS_969;
UNWINDOWED_970 <= FROM_DATAPATHS_970;
UNWINDOWED_971 <= FROM_DATAPATHS_971;
UNWINDOWED_972 <= FROM_DATAPATHS_972;
UNWINDOWED_973 <= FROM_DATAPATHS_973;
UNWINDOWED_974 <= FROM_DATAPATHS_974;
UNWINDOWED_975 <= FROM_DATAPATHS_975;
UNWINDOWED_976 <= FROM_DATAPATHS_976;
UNWINDOWED_977 <= FROM_DATAPATHS_977;
UNWINDOWED_978 <= FROM_DATAPATHS_978;
UNWINDOWED_979 <= FROM_DATAPATHS_979;
UNWINDOWED_980 <= FROM_DATAPATHS_980;
UNWINDOWED_981 <= FROM_DATAPATHS_981;
UNWINDOWED_982 <= FROM_DATAPATHS_982;
UNWINDOWED_983 <= FROM_DATAPATHS_983;
UNWINDOWED_984 <= FROM_DATAPATHS_984;
UNWINDOWED_985 <= FROM_DATAPATHS_985;
UNWINDOWED_986 <= FROM_DATAPATHS_986;
UNWINDOWED_987 <= FROM_DATAPATHS_987;
UNWINDOWED_988 <= FROM_DATAPATHS_988;
UNWINDOWED_989 <= FROM_DATAPATHS_989;
UNWINDOWED_990 <= FROM_DATAPATHS_990;
UNWINDOWED_991 <= FROM_DATAPATHS_991;
UNWINDOWED_992 <= FROM_DATAPATHS_992;
UNWINDOWED_993 <= FROM_DATAPATHS_993;
UNWINDOWED_994 <= FROM_DATAPATHS_994;
UNWINDOWED_995 <= FROM_DATAPATHS_995;
UNWINDOWED_996 <= FROM_DATAPATHS_996;
UNWINDOWED_997 <= FROM_DATAPATHS_997;
UNWINDOWED_998 <= FROM_DATAPATHS_998;
UNWINDOWED_999 <= FROM_DATAPATHS_999;
UNWINDOWED_1000 <= FROM_DATAPATHS_1000;
UNWINDOWED_1001 <= FROM_DATAPATHS_1001;
UNWINDOWED_1002 <= FROM_DATAPATHS_1002;
UNWINDOWED_1003 <= FROM_DATAPATHS_1003;
UNWINDOWED_1004 <= FROM_DATAPATHS_1004;
UNWINDOWED_1005 <= FROM_DATAPATHS_1005;
UNWINDOWED_1006 <= FROM_DATAPATHS_1006;
UNWINDOWED_1007 <= FROM_DATAPATHS_1007;
UNWINDOWED_1008 <= FROM_DATAPATHS_1008;
UNWINDOWED_1009 <= FROM_DATAPATHS_1009;
UNWINDOWED_1010 <= FROM_DATAPATHS_1010;
UNWINDOWED_1011 <= FROM_DATAPATHS_1011;
UNWINDOWED_1012 <= FROM_DATAPATHS_1012;
UNWINDOWED_1013 <= FROM_DATAPATHS_1013;
UNWINDOWED_1014 <= FROM_DATAPATHS_1014;
UNWINDOWED_1015 <= FROM_DATAPATHS_1015;
UNWINDOWED_1016 <= FROM_DATAPATHS_1016;
UNWINDOWED_1017 <= FROM_DATAPATHS_1017;
UNWINDOWED_1018 <= FROM_DATAPATHS_1018;
UNWINDOWED_1019 <= FROM_DATAPATHS_1019;
UNWINDOWED_1020 <= FROM_DATAPATHS_1020;
UNWINDOWED_1021 <= FROM_DATAPATHS_1021;
UNWINDOWED_1022 <= FROM_DATAPATHS_1022;
UNWINDOWED_1023 <= FROM_DATAPATHS_1023;

MUX_REORD_UNIT_0 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_0 ,
										MUX_10_1_IN_1 => UNWINDOWED_0 ,
										MUX_10_1_IN_2 => UNWINDOWED_0 ,
										MUX_10_1_IN_3 => UNWINDOWED_0 ,
										MUX_10_1_IN_4 => UNWINDOWED_0 ,
										MUX_10_1_IN_5 => UNWINDOWED_0 ,
										MUX_10_1_IN_6 => UNWINDOWED_0 ,
										MUX_10_1_IN_7 => UNWINDOWED_0 ,
										MUX_10_1_IN_8 => UNWINDOWED_0 ,
										MUX_10_1_IN_9 => UNWINDOWED_0 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_0
									);
MUX_REORD_UNIT_1 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1 ,
										MUX_10_1_IN_1 => UNWINDOWED_2 ,
										MUX_10_1_IN_2 => UNWINDOWED_2 ,
										MUX_10_1_IN_3 => UNWINDOWED_2 ,
										MUX_10_1_IN_4 => UNWINDOWED_2 ,
										MUX_10_1_IN_5 => UNWINDOWED_2 ,
										MUX_10_1_IN_6 => UNWINDOWED_2 ,
										MUX_10_1_IN_7 => UNWINDOWED_2 ,
										MUX_10_1_IN_8 => UNWINDOWED_2 ,
										MUX_10_1_IN_9 => UNWINDOWED_2 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1
									);
MUX_REORD_UNIT_2 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_2 ,
										MUX_10_1_IN_1 => UNWINDOWED_1 ,
										MUX_10_1_IN_2 => UNWINDOWED_4 ,
										MUX_10_1_IN_3 => UNWINDOWED_4 ,
										MUX_10_1_IN_4 => UNWINDOWED_4 ,
										MUX_10_1_IN_5 => UNWINDOWED_4 ,
										MUX_10_1_IN_6 => UNWINDOWED_4 ,
										MUX_10_1_IN_7 => UNWINDOWED_4 ,
										MUX_10_1_IN_8 => UNWINDOWED_4 ,
										MUX_10_1_IN_9 => UNWINDOWED_4 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_2
									);
MUX_REORD_UNIT_3 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_3 ,
										MUX_10_1_IN_1 => UNWINDOWED_3 ,
										MUX_10_1_IN_2 => UNWINDOWED_6 ,
										MUX_10_1_IN_3 => UNWINDOWED_6 ,
										MUX_10_1_IN_4 => UNWINDOWED_6 ,
										MUX_10_1_IN_5 => UNWINDOWED_6 ,
										MUX_10_1_IN_6 => UNWINDOWED_6 ,
										MUX_10_1_IN_7 => UNWINDOWED_6 ,
										MUX_10_1_IN_8 => UNWINDOWED_6 ,
										MUX_10_1_IN_9 => UNWINDOWED_6 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_3
									);
MUX_REORD_UNIT_4 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_4 ,
										MUX_10_1_IN_1 => UNWINDOWED_4 ,
										MUX_10_1_IN_2 => UNWINDOWED_1 ,
										MUX_10_1_IN_3 => UNWINDOWED_8 ,
										MUX_10_1_IN_4 => UNWINDOWED_8 ,
										MUX_10_1_IN_5 => UNWINDOWED_8 ,
										MUX_10_1_IN_6 => UNWINDOWED_8 ,
										MUX_10_1_IN_7 => UNWINDOWED_8 ,
										MUX_10_1_IN_8 => UNWINDOWED_8 ,
										MUX_10_1_IN_9 => UNWINDOWED_8 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_4
									);
MUX_REORD_UNIT_5 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_5 ,
										MUX_10_1_IN_1 => UNWINDOWED_6 ,
										MUX_10_1_IN_2 => UNWINDOWED_3 ,
										MUX_10_1_IN_3 => UNWINDOWED_10 ,
										MUX_10_1_IN_4 => UNWINDOWED_10 ,
										MUX_10_1_IN_5 => UNWINDOWED_10 ,
										MUX_10_1_IN_6 => UNWINDOWED_10 ,
										MUX_10_1_IN_7 => UNWINDOWED_10 ,
										MUX_10_1_IN_8 => UNWINDOWED_10 ,
										MUX_10_1_IN_9 => UNWINDOWED_10 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_5
									);
MUX_REORD_UNIT_6 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_6 ,
										MUX_10_1_IN_1 => UNWINDOWED_5 ,
										MUX_10_1_IN_2 => UNWINDOWED_5 ,
										MUX_10_1_IN_3 => UNWINDOWED_12 ,
										MUX_10_1_IN_4 => UNWINDOWED_12 ,
										MUX_10_1_IN_5 => UNWINDOWED_12 ,
										MUX_10_1_IN_6 => UNWINDOWED_12 ,
										MUX_10_1_IN_7 => UNWINDOWED_12 ,
										MUX_10_1_IN_8 => UNWINDOWED_12 ,
										MUX_10_1_IN_9 => UNWINDOWED_12 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_6
									);
MUX_REORD_UNIT_7 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_7 ,
										MUX_10_1_IN_1 => UNWINDOWED_7 ,
										MUX_10_1_IN_2 => UNWINDOWED_7 ,
										MUX_10_1_IN_3 => UNWINDOWED_14 ,
										MUX_10_1_IN_4 => UNWINDOWED_14 ,
										MUX_10_1_IN_5 => UNWINDOWED_14 ,
										MUX_10_1_IN_6 => UNWINDOWED_14 ,
										MUX_10_1_IN_7 => UNWINDOWED_14 ,
										MUX_10_1_IN_8 => UNWINDOWED_14 ,
										MUX_10_1_IN_9 => UNWINDOWED_14 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_7
									);
MUX_REORD_UNIT_8 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_8 ,
										MUX_10_1_IN_1 => UNWINDOWED_8 ,
										MUX_10_1_IN_2 => UNWINDOWED_8 ,
										MUX_10_1_IN_3 => UNWINDOWED_1 ,
										MUX_10_1_IN_4 => UNWINDOWED_16 ,
										MUX_10_1_IN_5 => UNWINDOWED_16 ,
										MUX_10_1_IN_6 => UNWINDOWED_16 ,
										MUX_10_1_IN_7 => UNWINDOWED_16 ,
										MUX_10_1_IN_8 => UNWINDOWED_16 ,
										MUX_10_1_IN_9 => UNWINDOWED_16 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_8
									);
MUX_REORD_UNIT_9 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_9 ,
										MUX_10_1_IN_1 => UNWINDOWED_10 ,
										MUX_10_1_IN_2 => UNWINDOWED_10 ,
										MUX_10_1_IN_3 => UNWINDOWED_3 ,
										MUX_10_1_IN_4 => UNWINDOWED_18 ,
										MUX_10_1_IN_5 => UNWINDOWED_18 ,
										MUX_10_1_IN_6 => UNWINDOWED_18 ,
										MUX_10_1_IN_7 => UNWINDOWED_18 ,
										MUX_10_1_IN_8 => UNWINDOWED_18 ,
										MUX_10_1_IN_9 => UNWINDOWED_18 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_9
									);
MUX_REORD_UNIT_10 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_10 ,
										MUX_10_1_IN_1 => UNWINDOWED_9 ,
										MUX_10_1_IN_2 => UNWINDOWED_12 ,
										MUX_10_1_IN_3 => UNWINDOWED_5 ,
										MUX_10_1_IN_4 => UNWINDOWED_20 ,
										MUX_10_1_IN_5 => UNWINDOWED_20 ,
										MUX_10_1_IN_6 => UNWINDOWED_20 ,
										MUX_10_1_IN_7 => UNWINDOWED_20 ,
										MUX_10_1_IN_8 => UNWINDOWED_20 ,
										MUX_10_1_IN_9 => UNWINDOWED_20 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_10
									);
MUX_REORD_UNIT_11 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_11 ,
										MUX_10_1_IN_1 => UNWINDOWED_11 ,
										MUX_10_1_IN_2 => UNWINDOWED_14 ,
										MUX_10_1_IN_3 => UNWINDOWED_7 ,
										MUX_10_1_IN_4 => UNWINDOWED_22 ,
										MUX_10_1_IN_5 => UNWINDOWED_22 ,
										MUX_10_1_IN_6 => UNWINDOWED_22 ,
										MUX_10_1_IN_7 => UNWINDOWED_22 ,
										MUX_10_1_IN_8 => UNWINDOWED_22 ,
										MUX_10_1_IN_9 => UNWINDOWED_22 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_11
									);
MUX_REORD_UNIT_12 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_12 ,
										MUX_10_1_IN_1 => UNWINDOWED_12 ,
										MUX_10_1_IN_2 => UNWINDOWED_9 ,
										MUX_10_1_IN_3 => UNWINDOWED_9 ,
										MUX_10_1_IN_4 => UNWINDOWED_24 ,
										MUX_10_1_IN_5 => UNWINDOWED_24 ,
										MUX_10_1_IN_6 => UNWINDOWED_24 ,
										MUX_10_1_IN_7 => UNWINDOWED_24 ,
										MUX_10_1_IN_8 => UNWINDOWED_24 ,
										MUX_10_1_IN_9 => UNWINDOWED_24 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_12
									);
MUX_REORD_UNIT_13 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_13 ,
										MUX_10_1_IN_1 => UNWINDOWED_14 ,
										MUX_10_1_IN_2 => UNWINDOWED_11 ,
										MUX_10_1_IN_3 => UNWINDOWED_11 ,
										MUX_10_1_IN_4 => UNWINDOWED_26 ,
										MUX_10_1_IN_5 => UNWINDOWED_26 ,
										MUX_10_1_IN_6 => UNWINDOWED_26 ,
										MUX_10_1_IN_7 => UNWINDOWED_26 ,
										MUX_10_1_IN_8 => UNWINDOWED_26 ,
										MUX_10_1_IN_9 => UNWINDOWED_26 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_13
									);
MUX_REORD_UNIT_14 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_14 ,
										MUX_10_1_IN_1 => UNWINDOWED_13 ,
										MUX_10_1_IN_2 => UNWINDOWED_13 ,
										MUX_10_1_IN_3 => UNWINDOWED_13 ,
										MUX_10_1_IN_4 => UNWINDOWED_28 ,
										MUX_10_1_IN_5 => UNWINDOWED_28 ,
										MUX_10_1_IN_6 => UNWINDOWED_28 ,
										MUX_10_1_IN_7 => UNWINDOWED_28 ,
										MUX_10_1_IN_8 => UNWINDOWED_28 ,
										MUX_10_1_IN_9 => UNWINDOWED_28 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_14
									);
MUX_REORD_UNIT_15 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_15 ,
										MUX_10_1_IN_1 => UNWINDOWED_15 ,
										MUX_10_1_IN_2 => UNWINDOWED_15 ,
										MUX_10_1_IN_3 => UNWINDOWED_15 ,
										MUX_10_1_IN_4 => UNWINDOWED_30 ,
										MUX_10_1_IN_5 => UNWINDOWED_30 ,
										MUX_10_1_IN_6 => UNWINDOWED_30 ,
										MUX_10_1_IN_7 => UNWINDOWED_30 ,
										MUX_10_1_IN_8 => UNWINDOWED_30 ,
										MUX_10_1_IN_9 => UNWINDOWED_30 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_15
									);
MUX_REORD_UNIT_16 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_16 ,
										MUX_10_1_IN_1 => UNWINDOWED_16 ,
										MUX_10_1_IN_2 => UNWINDOWED_16 ,
										MUX_10_1_IN_3 => UNWINDOWED_16 ,
										MUX_10_1_IN_4 => UNWINDOWED_1 ,
										MUX_10_1_IN_5 => UNWINDOWED_32 ,
										MUX_10_1_IN_6 => UNWINDOWED_32 ,
										MUX_10_1_IN_7 => UNWINDOWED_32 ,
										MUX_10_1_IN_8 => UNWINDOWED_32 ,
										MUX_10_1_IN_9 => UNWINDOWED_32 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_16
									);
MUX_REORD_UNIT_17 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_17 ,
										MUX_10_1_IN_1 => UNWINDOWED_18 ,
										MUX_10_1_IN_2 => UNWINDOWED_18 ,
										MUX_10_1_IN_3 => UNWINDOWED_18 ,
										MUX_10_1_IN_4 => UNWINDOWED_3 ,
										MUX_10_1_IN_5 => UNWINDOWED_34 ,
										MUX_10_1_IN_6 => UNWINDOWED_34 ,
										MUX_10_1_IN_7 => UNWINDOWED_34 ,
										MUX_10_1_IN_8 => UNWINDOWED_34 ,
										MUX_10_1_IN_9 => UNWINDOWED_34 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_17
									);
MUX_REORD_UNIT_18 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_18 ,
										MUX_10_1_IN_1 => UNWINDOWED_17 ,
										MUX_10_1_IN_2 => UNWINDOWED_20 ,
										MUX_10_1_IN_3 => UNWINDOWED_20 ,
										MUX_10_1_IN_4 => UNWINDOWED_5 ,
										MUX_10_1_IN_5 => UNWINDOWED_36 ,
										MUX_10_1_IN_6 => UNWINDOWED_36 ,
										MUX_10_1_IN_7 => UNWINDOWED_36 ,
										MUX_10_1_IN_8 => UNWINDOWED_36 ,
										MUX_10_1_IN_9 => UNWINDOWED_36 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_18
									);
MUX_REORD_UNIT_19 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_19 ,
										MUX_10_1_IN_1 => UNWINDOWED_19 ,
										MUX_10_1_IN_2 => UNWINDOWED_22 ,
										MUX_10_1_IN_3 => UNWINDOWED_22 ,
										MUX_10_1_IN_4 => UNWINDOWED_7 ,
										MUX_10_1_IN_5 => UNWINDOWED_38 ,
										MUX_10_1_IN_6 => UNWINDOWED_38 ,
										MUX_10_1_IN_7 => UNWINDOWED_38 ,
										MUX_10_1_IN_8 => UNWINDOWED_38 ,
										MUX_10_1_IN_9 => UNWINDOWED_38 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_19
									);
MUX_REORD_UNIT_20 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_20 ,
										MUX_10_1_IN_1 => UNWINDOWED_20 ,
										MUX_10_1_IN_2 => UNWINDOWED_17 ,
										MUX_10_1_IN_3 => UNWINDOWED_24 ,
										MUX_10_1_IN_4 => UNWINDOWED_9 ,
										MUX_10_1_IN_5 => UNWINDOWED_40 ,
										MUX_10_1_IN_6 => UNWINDOWED_40 ,
										MUX_10_1_IN_7 => UNWINDOWED_40 ,
										MUX_10_1_IN_8 => UNWINDOWED_40 ,
										MUX_10_1_IN_9 => UNWINDOWED_40 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_20
									);
MUX_REORD_UNIT_21 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_21 ,
										MUX_10_1_IN_1 => UNWINDOWED_22 ,
										MUX_10_1_IN_2 => UNWINDOWED_19 ,
										MUX_10_1_IN_3 => UNWINDOWED_26 ,
										MUX_10_1_IN_4 => UNWINDOWED_11 ,
										MUX_10_1_IN_5 => UNWINDOWED_42 ,
										MUX_10_1_IN_6 => UNWINDOWED_42 ,
										MUX_10_1_IN_7 => UNWINDOWED_42 ,
										MUX_10_1_IN_8 => UNWINDOWED_42 ,
										MUX_10_1_IN_9 => UNWINDOWED_42 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_21
									);
MUX_REORD_UNIT_22 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_22 ,
										MUX_10_1_IN_1 => UNWINDOWED_21 ,
										MUX_10_1_IN_2 => UNWINDOWED_21 ,
										MUX_10_1_IN_3 => UNWINDOWED_28 ,
										MUX_10_1_IN_4 => UNWINDOWED_13 ,
										MUX_10_1_IN_5 => UNWINDOWED_44 ,
										MUX_10_1_IN_6 => UNWINDOWED_44 ,
										MUX_10_1_IN_7 => UNWINDOWED_44 ,
										MUX_10_1_IN_8 => UNWINDOWED_44 ,
										MUX_10_1_IN_9 => UNWINDOWED_44 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_22
									);
MUX_REORD_UNIT_23 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_23 ,
										MUX_10_1_IN_1 => UNWINDOWED_23 ,
										MUX_10_1_IN_2 => UNWINDOWED_23 ,
										MUX_10_1_IN_3 => UNWINDOWED_30 ,
										MUX_10_1_IN_4 => UNWINDOWED_15 ,
										MUX_10_1_IN_5 => UNWINDOWED_46 ,
										MUX_10_1_IN_6 => UNWINDOWED_46 ,
										MUX_10_1_IN_7 => UNWINDOWED_46 ,
										MUX_10_1_IN_8 => UNWINDOWED_46 ,
										MUX_10_1_IN_9 => UNWINDOWED_46 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_23
									);
MUX_REORD_UNIT_24 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_24 ,
										MUX_10_1_IN_1 => UNWINDOWED_24 ,
										MUX_10_1_IN_2 => UNWINDOWED_24 ,
										MUX_10_1_IN_3 => UNWINDOWED_17 ,
										MUX_10_1_IN_4 => UNWINDOWED_17 ,
										MUX_10_1_IN_5 => UNWINDOWED_48 ,
										MUX_10_1_IN_6 => UNWINDOWED_48 ,
										MUX_10_1_IN_7 => UNWINDOWED_48 ,
										MUX_10_1_IN_8 => UNWINDOWED_48 ,
										MUX_10_1_IN_9 => UNWINDOWED_48 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_24
									);
MUX_REORD_UNIT_25 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_25 ,
										MUX_10_1_IN_1 => UNWINDOWED_26 ,
										MUX_10_1_IN_2 => UNWINDOWED_26 ,
										MUX_10_1_IN_3 => UNWINDOWED_19 ,
										MUX_10_1_IN_4 => UNWINDOWED_19 ,
										MUX_10_1_IN_5 => UNWINDOWED_50 ,
										MUX_10_1_IN_6 => UNWINDOWED_50 ,
										MUX_10_1_IN_7 => UNWINDOWED_50 ,
										MUX_10_1_IN_8 => UNWINDOWED_50 ,
										MUX_10_1_IN_9 => UNWINDOWED_50 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_25
									);
MUX_REORD_UNIT_26 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_26 ,
										MUX_10_1_IN_1 => UNWINDOWED_25 ,
										MUX_10_1_IN_2 => UNWINDOWED_28 ,
										MUX_10_1_IN_3 => UNWINDOWED_21 ,
										MUX_10_1_IN_4 => UNWINDOWED_21 ,
										MUX_10_1_IN_5 => UNWINDOWED_52 ,
										MUX_10_1_IN_6 => UNWINDOWED_52 ,
										MUX_10_1_IN_7 => UNWINDOWED_52 ,
										MUX_10_1_IN_8 => UNWINDOWED_52 ,
										MUX_10_1_IN_9 => UNWINDOWED_52 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_26
									);
MUX_REORD_UNIT_27 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_27 ,
										MUX_10_1_IN_1 => UNWINDOWED_27 ,
										MUX_10_1_IN_2 => UNWINDOWED_30 ,
										MUX_10_1_IN_3 => UNWINDOWED_23 ,
										MUX_10_1_IN_4 => UNWINDOWED_23 ,
										MUX_10_1_IN_5 => UNWINDOWED_54 ,
										MUX_10_1_IN_6 => UNWINDOWED_54 ,
										MUX_10_1_IN_7 => UNWINDOWED_54 ,
										MUX_10_1_IN_8 => UNWINDOWED_54 ,
										MUX_10_1_IN_9 => UNWINDOWED_54 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_27
									);
MUX_REORD_UNIT_28 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_28 ,
										MUX_10_1_IN_1 => UNWINDOWED_28 ,
										MUX_10_1_IN_2 => UNWINDOWED_25 ,
										MUX_10_1_IN_3 => UNWINDOWED_25 ,
										MUX_10_1_IN_4 => UNWINDOWED_25 ,
										MUX_10_1_IN_5 => UNWINDOWED_56 ,
										MUX_10_1_IN_6 => UNWINDOWED_56 ,
										MUX_10_1_IN_7 => UNWINDOWED_56 ,
										MUX_10_1_IN_8 => UNWINDOWED_56 ,
										MUX_10_1_IN_9 => UNWINDOWED_56 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_28
									);
MUX_REORD_UNIT_29 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_29 ,
										MUX_10_1_IN_1 => UNWINDOWED_30 ,
										MUX_10_1_IN_2 => UNWINDOWED_27 ,
										MUX_10_1_IN_3 => UNWINDOWED_27 ,
										MUX_10_1_IN_4 => UNWINDOWED_27 ,
										MUX_10_1_IN_5 => UNWINDOWED_58 ,
										MUX_10_1_IN_6 => UNWINDOWED_58 ,
										MUX_10_1_IN_7 => UNWINDOWED_58 ,
										MUX_10_1_IN_8 => UNWINDOWED_58 ,
										MUX_10_1_IN_9 => UNWINDOWED_58 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_29
									);
MUX_REORD_UNIT_30 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_30 ,
										MUX_10_1_IN_1 => UNWINDOWED_29 ,
										MUX_10_1_IN_2 => UNWINDOWED_29 ,
										MUX_10_1_IN_3 => UNWINDOWED_29 ,
										MUX_10_1_IN_4 => UNWINDOWED_29 ,
										MUX_10_1_IN_5 => UNWINDOWED_60 ,
										MUX_10_1_IN_6 => UNWINDOWED_60 ,
										MUX_10_1_IN_7 => UNWINDOWED_60 ,
										MUX_10_1_IN_8 => UNWINDOWED_60 ,
										MUX_10_1_IN_9 => UNWINDOWED_60 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_30
									);
MUX_REORD_UNIT_31 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_31 ,
										MUX_10_1_IN_1 => UNWINDOWED_31 ,
										MUX_10_1_IN_2 => UNWINDOWED_31 ,
										MUX_10_1_IN_3 => UNWINDOWED_31 ,
										MUX_10_1_IN_4 => UNWINDOWED_31 ,
										MUX_10_1_IN_5 => UNWINDOWED_62 ,
										MUX_10_1_IN_6 => UNWINDOWED_62 ,
										MUX_10_1_IN_7 => UNWINDOWED_62 ,
										MUX_10_1_IN_8 => UNWINDOWED_62 ,
										MUX_10_1_IN_9 => UNWINDOWED_62 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_31
									);
MUX_REORD_UNIT_32 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_32 ,
										MUX_10_1_IN_1 => UNWINDOWED_32 ,
										MUX_10_1_IN_2 => UNWINDOWED_32 ,
										MUX_10_1_IN_3 => UNWINDOWED_32 ,
										MUX_10_1_IN_4 => UNWINDOWED_32 ,
										MUX_10_1_IN_5 => UNWINDOWED_1 ,
										MUX_10_1_IN_6 => UNWINDOWED_64 ,
										MUX_10_1_IN_7 => UNWINDOWED_64 ,
										MUX_10_1_IN_8 => UNWINDOWED_64 ,
										MUX_10_1_IN_9 => UNWINDOWED_64 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_32
									);
MUX_REORD_UNIT_33 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_33 ,
										MUX_10_1_IN_1 => UNWINDOWED_34 ,
										MUX_10_1_IN_2 => UNWINDOWED_34 ,
										MUX_10_1_IN_3 => UNWINDOWED_34 ,
										MUX_10_1_IN_4 => UNWINDOWED_34 ,
										MUX_10_1_IN_5 => UNWINDOWED_3 ,
										MUX_10_1_IN_6 => UNWINDOWED_66 ,
										MUX_10_1_IN_7 => UNWINDOWED_66 ,
										MUX_10_1_IN_8 => UNWINDOWED_66 ,
										MUX_10_1_IN_9 => UNWINDOWED_66 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_33
									);
MUX_REORD_UNIT_34 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_34 ,
										MUX_10_1_IN_1 => UNWINDOWED_33 ,
										MUX_10_1_IN_2 => UNWINDOWED_36 ,
										MUX_10_1_IN_3 => UNWINDOWED_36 ,
										MUX_10_1_IN_4 => UNWINDOWED_36 ,
										MUX_10_1_IN_5 => UNWINDOWED_5 ,
										MUX_10_1_IN_6 => UNWINDOWED_68 ,
										MUX_10_1_IN_7 => UNWINDOWED_68 ,
										MUX_10_1_IN_8 => UNWINDOWED_68 ,
										MUX_10_1_IN_9 => UNWINDOWED_68 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_34
									);
MUX_REORD_UNIT_35 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_35 ,
										MUX_10_1_IN_1 => UNWINDOWED_35 ,
										MUX_10_1_IN_2 => UNWINDOWED_38 ,
										MUX_10_1_IN_3 => UNWINDOWED_38 ,
										MUX_10_1_IN_4 => UNWINDOWED_38 ,
										MUX_10_1_IN_5 => UNWINDOWED_7 ,
										MUX_10_1_IN_6 => UNWINDOWED_70 ,
										MUX_10_1_IN_7 => UNWINDOWED_70 ,
										MUX_10_1_IN_8 => UNWINDOWED_70 ,
										MUX_10_1_IN_9 => UNWINDOWED_70 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_35
									);
MUX_REORD_UNIT_36 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_36 ,
										MUX_10_1_IN_1 => UNWINDOWED_36 ,
										MUX_10_1_IN_2 => UNWINDOWED_33 ,
										MUX_10_1_IN_3 => UNWINDOWED_40 ,
										MUX_10_1_IN_4 => UNWINDOWED_40 ,
										MUX_10_1_IN_5 => UNWINDOWED_9 ,
										MUX_10_1_IN_6 => UNWINDOWED_72 ,
										MUX_10_1_IN_7 => UNWINDOWED_72 ,
										MUX_10_1_IN_8 => UNWINDOWED_72 ,
										MUX_10_1_IN_9 => UNWINDOWED_72 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_36
									);
MUX_REORD_UNIT_37 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_37 ,
										MUX_10_1_IN_1 => UNWINDOWED_38 ,
										MUX_10_1_IN_2 => UNWINDOWED_35 ,
										MUX_10_1_IN_3 => UNWINDOWED_42 ,
										MUX_10_1_IN_4 => UNWINDOWED_42 ,
										MUX_10_1_IN_5 => UNWINDOWED_11 ,
										MUX_10_1_IN_6 => UNWINDOWED_74 ,
										MUX_10_1_IN_7 => UNWINDOWED_74 ,
										MUX_10_1_IN_8 => UNWINDOWED_74 ,
										MUX_10_1_IN_9 => UNWINDOWED_74 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_37
									);
MUX_REORD_UNIT_38 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_38 ,
										MUX_10_1_IN_1 => UNWINDOWED_37 ,
										MUX_10_1_IN_2 => UNWINDOWED_37 ,
										MUX_10_1_IN_3 => UNWINDOWED_44 ,
										MUX_10_1_IN_4 => UNWINDOWED_44 ,
										MUX_10_1_IN_5 => UNWINDOWED_13 ,
										MUX_10_1_IN_6 => UNWINDOWED_76 ,
										MUX_10_1_IN_7 => UNWINDOWED_76 ,
										MUX_10_1_IN_8 => UNWINDOWED_76 ,
										MUX_10_1_IN_9 => UNWINDOWED_76 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_38
									);
MUX_REORD_UNIT_39 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_39 ,
										MUX_10_1_IN_1 => UNWINDOWED_39 ,
										MUX_10_1_IN_2 => UNWINDOWED_39 ,
										MUX_10_1_IN_3 => UNWINDOWED_46 ,
										MUX_10_1_IN_4 => UNWINDOWED_46 ,
										MUX_10_1_IN_5 => UNWINDOWED_15 ,
										MUX_10_1_IN_6 => UNWINDOWED_78 ,
										MUX_10_1_IN_7 => UNWINDOWED_78 ,
										MUX_10_1_IN_8 => UNWINDOWED_78 ,
										MUX_10_1_IN_9 => UNWINDOWED_78 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_39
									);
MUX_REORD_UNIT_40 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_40 ,
										MUX_10_1_IN_1 => UNWINDOWED_40 ,
										MUX_10_1_IN_2 => UNWINDOWED_40 ,
										MUX_10_1_IN_3 => UNWINDOWED_33 ,
										MUX_10_1_IN_4 => UNWINDOWED_48 ,
										MUX_10_1_IN_5 => UNWINDOWED_17 ,
										MUX_10_1_IN_6 => UNWINDOWED_80 ,
										MUX_10_1_IN_7 => UNWINDOWED_80 ,
										MUX_10_1_IN_8 => UNWINDOWED_80 ,
										MUX_10_1_IN_9 => UNWINDOWED_80 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_40
									);
MUX_REORD_UNIT_41 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_41 ,
										MUX_10_1_IN_1 => UNWINDOWED_42 ,
										MUX_10_1_IN_2 => UNWINDOWED_42 ,
										MUX_10_1_IN_3 => UNWINDOWED_35 ,
										MUX_10_1_IN_4 => UNWINDOWED_50 ,
										MUX_10_1_IN_5 => UNWINDOWED_19 ,
										MUX_10_1_IN_6 => UNWINDOWED_82 ,
										MUX_10_1_IN_7 => UNWINDOWED_82 ,
										MUX_10_1_IN_8 => UNWINDOWED_82 ,
										MUX_10_1_IN_9 => UNWINDOWED_82 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_41
									);
MUX_REORD_UNIT_42 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_42 ,
										MUX_10_1_IN_1 => UNWINDOWED_41 ,
										MUX_10_1_IN_2 => UNWINDOWED_44 ,
										MUX_10_1_IN_3 => UNWINDOWED_37 ,
										MUX_10_1_IN_4 => UNWINDOWED_52 ,
										MUX_10_1_IN_5 => UNWINDOWED_21 ,
										MUX_10_1_IN_6 => UNWINDOWED_84 ,
										MUX_10_1_IN_7 => UNWINDOWED_84 ,
										MUX_10_1_IN_8 => UNWINDOWED_84 ,
										MUX_10_1_IN_9 => UNWINDOWED_84 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_42
									);
MUX_REORD_UNIT_43 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_43 ,
										MUX_10_1_IN_1 => UNWINDOWED_43 ,
										MUX_10_1_IN_2 => UNWINDOWED_46 ,
										MUX_10_1_IN_3 => UNWINDOWED_39 ,
										MUX_10_1_IN_4 => UNWINDOWED_54 ,
										MUX_10_1_IN_5 => UNWINDOWED_23 ,
										MUX_10_1_IN_6 => UNWINDOWED_86 ,
										MUX_10_1_IN_7 => UNWINDOWED_86 ,
										MUX_10_1_IN_8 => UNWINDOWED_86 ,
										MUX_10_1_IN_9 => UNWINDOWED_86 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_43
									);
MUX_REORD_UNIT_44 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_44 ,
										MUX_10_1_IN_1 => UNWINDOWED_44 ,
										MUX_10_1_IN_2 => UNWINDOWED_41 ,
										MUX_10_1_IN_3 => UNWINDOWED_41 ,
										MUX_10_1_IN_4 => UNWINDOWED_56 ,
										MUX_10_1_IN_5 => UNWINDOWED_25 ,
										MUX_10_1_IN_6 => UNWINDOWED_88 ,
										MUX_10_1_IN_7 => UNWINDOWED_88 ,
										MUX_10_1_IN_8 => UNWINDOWED_88 ,
										MUX_10_1_IN_9 => UNWINDOWED_88 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_44
									);
MUX_REORD_UNIT_45 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_45 ,
										MUX_10_1_IN_1 => UNWINDOWED_46 ,
										MUX_10_1_IN_2 => UNWINDOWED_43 ,
										MUX_10_1_IN_3 => UNWINDOWED_43 ,
										MUX_10_1_IN_4 => UNWINDOWED_58 ,
										MUX_10_1_IN_5 => UNWINDOWED_27 ,
										MUX_10_1_IN_6 => UNWINDOWED_90 ,
										MUX_10_1_IN_7 => UNWINDOWED_90 ,
										MUX_10_1_IN_8 => UNWINDOWED_90 ,
										MUX_10_1_IN_9 => UNWINDOWED_90 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_45
									);
MUX_REORD_UNIT_46 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_46 ,
										MUX_10_1_IN_1 => UNWINDOWED_45 ,
										MUX_10_1_IN_2 => UNWINDOWED_45 ,
										MUX_10_1_IN_3 => UNWINDOWED_45 ,
										MUX_10_1_IN_4 => UNWINDOWED_60 ,
										MUX_10_1_IN_5 => UNWINDOWED_29 ,
										MUX_10_1_IN_6 => UNWINDOWED_92 ,
										MUX_10_1_IN_7 => UNWINDOWED_92 ,
										MUX_10_1_IN_8 => UNWINDOWED_92 ,
										MUX_10_1_IN_9 => UNWINDOWED_92 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_46
									);
MUX_REORD_UNIT_47 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_47 ,
										MUX_10_1_IN_1 => UNWINDOWED_47 ,
										MUX_10_1_IN_2 => UNWINDOWED_47 ,
										MUX_10_1_IN_3 => UNWINDOWED_47 ,
										MUX_10_1_IN_4 => UNWINDOWED_62 ,
										MUX_10_1_IN_5 => UNWINDOWED_31 ,
										MUX_10_1_IN_6 => UNWINDOWED_94 ,
										MUX_10_1_IN_7 => UNWINDOWED_94 ,
										MUX_10_1_IN_8 => UNWINDOWED_94 ,
										MUX_10_1_IN_9 => UNWINDOWED_94 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_47
									);
MUX_REORD_UNIT_48 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_48 ,
										MUX_10_1_IN_1 => UNWINDOWED_48 ,
										MUX_10_1_IN_2 => UNWINDOWED_48 ,
										MUX_10_1_IN_3 => UNWINDOWED_48 ,
										MUX_10_1_IN_4 => UNWINDOWED_33 ,
										MUX_10_1_IN_5 => UNWINDOWED_33 ,
										MUX_10_1_IN_6 => UNWINDOWED_96 ,
										MUX_10_1_IN_7 => UNWINDOWED_96 ,
										MUX_10_1_IN_8 => UNWINDOWED_96 ,
										MUX_10_1_IN_9 => UNWINDOWED_96 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_48
									);
MUX_REORD_UNIT_49 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_49 ,
										MUX_10_1_IN_1 => UNWINDOWED_50 ,
										MUX_10_1_IN_2 => UNWINDOWED_50 ,
										MUX_10_1_IN_3 => UNWINDOWED_50 ,
										MUX_10_1_IN_4 => UNWINDOWED_35 ,
										MUX_10_1_IN_5 => UNWINDOWED_35 ,
										MUX_10_1_IN_6 => UNWINDOWED_98 ,
										MUX_10_1_IN_7 => UNWINDOWED_98 ,
										MUX_10_1_IN_8 => UNWINDOWED_98 ,
										MUX_10_1_IN_9 => UNWINDOWED_98 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_49
									);
MUX_REORD_UNIT_50 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_50 ,
										MUX_10_1_IN_1 => UNWINDOWED_49 ,
										MUX_10_1_IN_2 => UNWINDOWED_52 ,
										MUX_10_1_IN_3 => UNWINDOWED_52 ,
										MUX_10_1_IN_4 => UNWINDOWED_37 ,
										MUX_10_1_IN_5 => UNWINDOWED_37 ,
										MUX_10_1_IN_6 => UNWINDOWED_100 ,
										MUX_10_1_IN_7 => UNWINDOWED_100 ,
										MUX_10_1_IN_8 => UNWINDOWED_100 ,
										MUX_10_1_IN_9 => UNWINDOWED_100 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_50
									);
MUX_REORD_UNIT_51 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_51 ,
										MUX_10_1_IN_1 => UNWINDOWED_51 ,
										MUX_10_1_IN_2 => UNWINDOWED_54 ,
										MUX_10_1_IN_3 => UNWINDOWED_54 ,
										MUX_10_1_IN_4 => UNWINDOWED_39 ,
										MUX_10_1_IN_5 => UNWINDOWED_39 ,
										MUX_10_1_IN_6 => UNWINDOWED_102 ,
										MUX_10_1_IN_7 => UNWINDOWED_102 ,
										MUX_10_1_IN_8 => UNWINDOWED_102 ,
										MUX_10_1_IN_9 => UNWINDOWED_102 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_51
									);
MUX_REORD_UNIT_52 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_52 ,
										MUX_10_1_IN_1 => UNWINDOWED_52 ,
										MUX_10_1_IN_2 => UNWINDOWED_49 ,
										MUX_10_1_IN_3 => UNWINDOWED_56 ,
										MUX_10_1_IN_4 => UNWINDOWED_41 ,
										MUX_10_1_IN_5 => UNWINDOWED_41 ,
										MUX_10_1_IN_6 => UNWINDOWED_104 ,
										MUX_10_1_IN_7 => UNWINDOWED_104 ,
										MUX_10_1_IN_8 => UNWINDOWED_104 ,
										MUX_10_1_IN_9 => UNWINDOWED_104 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_52
									);
MUX_REORD_UNIT_53 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_53 ,
										MUX_10_1_IN_1 => UNWINDOWED_54 ,
										MUX_10_1_IN_2 => UNWINDOWED_51 ,
										MUX_10_1_IN_3 => UNWINDOWED_58 ,
										MUX_10_1_IN_4 => UNWINDOWED_43 ,
										MUX_10_1_IN_5 => UNWINDOWED_43 ,
										MUX_10_1_IN_6 => UNWINDOWED_106 ,
										MUX_10_1_IN_7 => UNWINDOWED_106 ,
										MUX_10_1_IN_8 => UNWINDOWED_106 ,
										MUX_10_1_IN_9 => UNWINDOWED_106 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_53
									);
MUX_REORD_UNIT_54 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_54 ,
										MUX_10_1_IN_1 => UNWINDOWED_53 ,
										MUX_10_1_IN_2 => UNWINDOWED_53 ,
										MUX_10_1_IN_3 => UNWINDOWED_60 ,
										MUX_10_1_IN_4 => UNWINDOWED_45 ,
										MUX_10_1_IN_5 => UNWINDOWED_45 ,
										MUX_10_1_IN_6 => UNWINDOWED_108 ,
										MUX_10_1_IN_7 => UNWINDOWED_108 ,
										MUX_10_1_IN_8 => UNWINDOWED_108 ,
										MUX_10_1_IN_9 => UNWINDOWED_108 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_54
									);
MUX_REORD_UNIT_55 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_55 ,
										MUX_10_1_IN_1 => UNWINDOWED_55 ,
										MUX_10_1_IN_2 => UNWINDOWED_55 ,
										MUX_10_1_IN_3 => UNWINDOWED_62 ,
										MUX_10_1_IN_4 => UNWINDOWED_47 ,
										MUX_10_1_IN_5 => UNWINDOWED_47 ,
										MUX_10_1_IN_6 => UNWINDOWED_110 ,
										MUX_10_1_IN_7 => UNWINDOWED_110 ,
										MUX_10_1_IN_8 => UNWINDOWED_110 ,
										MUX_10_1_IN_9 => UNWINDOWED_110 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_55
									);
MUX_REORD_UNIT_56 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_56 ,
										MUX_10_1_IN_1 => UNWINDOWED_56 ,
										MUX_10_1_IN_2 => UNWINDOWED_56 ,
										MUX_10_1_IN_3 => UNWINDOWED_49 ,
										MUX_10_1_IN_4 => UNWINDOWED_49 ,
										MUX_10_1_IN_5 => UNWINDOWED_49 ,
										MUX_10_1_IN_6 => UNWINDOWED_112 ,
										MUX_10_1_IN_7 => UNWINDOWED_112 ,
										MUX_10_1_IN_8 => UNWINDOWED_112 ,
										MUX_10_1_IN_9 => UNWINDOWED_112 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_56
									);
MUX_REORD_UNIT_57 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_57 ,
										MUX_10_1_IN_1 => UNWINDOWED_58 ,
										MUX_10_1_IN_2 => UNWINDOWED_58 ,
										MUX_10_1_IN_3 => UNWINDOWED_51 ,
										MUX_10_1_IN_4 => UNWINDOWED_51 ,
										MUX_10_1_IN_5 => UNWINDOWED_51 ,
										MUX_10_1_IN_6 => UNWINDOWED_114 ,
										MUX_10_1_IN_7 => UNWINDOWED_114 ,
										MUX_10_1_IN_8 => UNWINDOWED_114 ,
										MUX_10_1_IN_9 => UNWINDOWED_114 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_57
									);
MUX_REORD_UNIT_58 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_58 ,
										MUX_10_1_IN_1 => UNWINDOWED_57 ,
										MUX_10_1_IN_2 => UNWINDOWED_60 ,
										MUX_10_1_IN_3 => UNWINDOWED_53 ,
										MUX_10_1_IN_4 => UNWINDOWED_53 ,
										MUX_10_1_IN_5 => UNWINDOWED_53 ,
										MUX_10_1_IN_6 => UNWINDOWED_116 ,
										MUX_10_1_IN_7 => UNWINDOWED_116 ,
										MUX_10_1_IN_8 => UNWINDOWED_116 ,
										MUX_10_1_IN_9 => UNWINDOWED_116 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_58
									);
MUX_REORD_UNIT_59 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_59 ,
										MUX_10_1_IN_1 => UNWINDOWED_59 ,
										MUX_10_1_IN_2 => UNWINDOWED_62 ,
										MUX_10_1_IN_3 => UNWINDOWED_55 ,
										MUX_10_1_IN_4 => UNWINDOWED_55 ,
										MUX_10_1_IN_5 => UNWINDOWED_55 ,
										MUX_10_1_IN_6 => UNWINDOWED_118 ,
										MUX_10_1_IN_7 => UNWINDOWED_118 ,
										MUX_10_1_IN_8 => UNWINDOWED_118 ,
										MUX_10_1_IN_9 => UNWINDOWED_118 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_59
									);
MUX_REORD_UNIT_60 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_60 ,
										MUX_10_1_IN_1 => UNWINDOWED_60 ,
										MUX_10_1_IN_2 => UNWINDOWED_57 ,
										MUX_10_1_IN_3 => UNWINDOWED_57 ,
										MUX_10_1_IN_4 => UNWINDOWED_57 ,
										MUX_10_1_IN_5 => UNWINDOWED_57 ,
										MUX_10_1_IN_6 => UNWINDOWED_120 ,
										MUX_10_1_IN_7 => UNWINDOWED_120 ,
										MUX_10_1_IN_8 => UNWINDOWED_120 ,
										MUX_10_1_IN_9 => UNWINDOWED_120 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_60
									);
MUX_REORD_UNIT_61 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_61 ,
										MUX_10_1_IN_1 => UNWINDOWED_62 ,
										MUX_10_1_IN_2 => UNWINDOWED_59 ,
										MUX_10_1_IN_3 => UNWINDOWED_59 ,
										MUX_10_1_IN_4 => UNWINDOWED_59 ,
										MUX_10_1_IN_5 => UNWINDOWED_59 ,
										MUX_10_1_IN_6 => UNWINDOWED_122 ,
										MUX_10_1_IN_7 => UNWINDOWED_122 ,
										MUX_10_1_IN_8 => UNWINDOWED_122 ,
										MUX_10_1_IN_9 => UNWINDOWED_122 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_61
									);
MUX_REORD_UNIT_62 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_62 ,
										MUX_10_1_IN_1 => UNWINDOWED_61 ,
										MUX_10_1_IN_2 => UNWINDOWED_61 ,
										MUX_10_1_IN_3 => UNWINDOWED_61 ,
										MUX_10_1_IN_4 => UNWINDOWED_61 ,
										MUX_10_1_IN_5 => UNWINDOWED_61 ,
										MUX_10_1_IN_6 => UNWINDOWED_124 ,
										MUX_10_1_IN_7 => UNWINDOWED_124 ,
										MUX_10_1_IN_8 => UNWINDOWED_124 ,
										MUX_10_1_IN_9 => UNWINDOWED_124 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_62
									);
MUX_REORD_UNIT_63 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_63 ,
										MUX_10_1_IN_1 => UNWINDOWED_63 ,
										MUX_10_1_IN_2 => UNWINDOWED_63 ,
										MUX_10_1_IN_3 => UNWINDOWED_63 ,
										MUX_10_1_IN_4 => UNWINDOWED_63 ,
										MUX_10_1_IN_5 => UNWINDOWED_63 ,
										MUX_10_1_IN_6 => UNWINDOWED_126 ,
										MUX_10_1_IN_7 => UNWINDOWED_126 ,
										MUX_10_1_IN_8 => UNWINDOWED_126 ,
										MUX_10_1_IN_9 => UNWINDOWED_126 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_63
									);
MUX_REORD_UNIT_64 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_64 ,
										MUX_10_1_IN_1 => UNWINDOWED_64 ,
										MUX_10_1_IN_2 => UNWINDOWED_64 ,
										MUX_10_1_IN_3 => UNWINDOWED_64 ,
										MUX_10_1_IN_4 => UNWINDOWED_64 ,
										MUX_10_1_IN_5 => UNWINDOWED_64 ,
										MUX_10_1_IN_6 => UNWINDOWED_1 ,
										MUX_10_1_IN_7 => UNWINDOWED_128 ,
										MUX_10_1_IN_8 => UNWINDOWED_128 ,
										MUX_10_1_IN_9 => UNWINDOWED_128 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_64
									);
MUX_REORD_UNIT_65 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_65 ,
										MUX_10_1_IN_1 => UNWINDOWED_66 ,
										MUX_10_1_IN_2 => UNWINDOWED_66 ,
										MUX_10_1_IN_3 => UNWINDOWED_66 ,
										MUX_10_1_IN_4 => UNWINDOWED_66 ,
										MUX_10_1_IN_5 => UNWINDOWED_66 ,
										MUX_10_1_IN_6 => UNWINDOWED_3 ,
										MUX_10_1_IN_7 => UNWINDOWED_130 ,
										MUX_10_1_IN_8 => UNWINDOWED_130 ,
										MUX_10_1_IN_9 => UNWINDOWED_130 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_65
									);
MUX_REORD_UNIT_66 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_66 ,
										MUX_10_1_IN_1 => UNWINDOWED_65 ,
										MUX_10_1_IN_2 => UNWINDOWED_68 ,
										MUX_10_1_IN_3 => UNWINDOWED_68 ,
										MUX_10_1_IN_4 => UNWINDOWED_68 ,
										MUX_10_1_IN_5 => UNWINDOWED_68 ,
										MUX_10_1_IN_6 => UNWINDOWED_5 ,
										MUX_10_1_IN_7 => UNWINDOWED_132 ,
										MUX_10_1_IN_8 => UNWINDOWED_132 ,
										MUX_10_1_IN_9 => UNWINDOWED_132 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_66
									);
MUX_REORD_UNIT_67 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_67 ,
										MUX_10_1_IN_1 => UNWINDOWED_67 ,
										MUX_10_1_IN_2 => UNWINDOWED_70 ,
										MUX_10_1_IN_3 => UNWINDOWED_70 ,
										MUX_10_1_IN_4 => UNWINDOWED_70 ,
										MUX_10_1_IN_5 => UNWINDOWED_70 ,
										MUX_10_1_IN_6 => UNWINDOWED_7 ,
										MUX_10_1_IN_7 => UNWINDOWED_134 ,
										MUX_10_1_IN_8 => UNWINDOWED_134 ,
										MUX_10_1_IN_9 => UNWINDOWED_134 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_67
									);
MUX_REORD_UNIT_68 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_68 ,
										MUX_10_1_IN_1 => UNWINDOWED_68 ,
										MUX_10_1_IN_2 => UNWINDOWED_65 ,
										MUX_10_1_IN_3 => UNWINDOWED_72 ,
										MUX_10_1_IN_4 => UNWINDOWED_72 ,
										MUX_10_1_IN_5 => UNWINDOWED_72 ,
										MUX_10_1_IN_6 => UNWINDOWED_9 ,
										MUX_10_1_IN_7 => UNWINDOWED_136 ,
										MUX_10_1_IN_8 => UNWINDOWED_136 ,
										MUX_10_1_IN_9 => UNWINDOWED_136 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_68
									);
MUX_REORD_UNIT_69 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_69 ,
										MUX_10_1_IN_1 => UNWINDOWED_70 ,
										MUX_10_1_IN_2 => UNWINDOWED_67 ,
										MUX_10_1_IN_3 => UNWINDOWED_74 ,
										MUX_10_1_IN_4 => UNWINDOWED_74 ,
										MUX_10_1_IN_5 => UNWINDOWED_74 ,
										MUX_10_1_IN_6 => UNWINDOWED_11 ,
										MUX_10_1_IN_7 => UNWINDOWED_138 ,
										MUX_10_1_IN_8 => UNWINDOWED_138 ,
										MUX_10_1_IN_9 => UNWINDOWED_138 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_69
									);
MUX_REORD_UNIT_70 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_70 ,
										MUX_10_1_IN_1 => UNWINDOWED_69 ,
										MUX_10_1_IN_2 => UNWINDOWED_69 ,
										MUX_10_1_IN_3 => UNWINDOWED_76 ,
										MUX_10_1_IN_4 => UNWINDOWED_76 ,
										MUX_10_1_IN_5 => UNWINDOWED_76 ,
										MUX_10_1_IN_6 => UNWINDOWED_13 ,
										MUX_10_1_IN_7 => UNWINDOWED_140 ,
										MUX_10_1_IN_8 => UNWINDOWED_140 ,
										MUX_10_1_IN_9 => UNWINDOWED_140 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_70
									);
MUX_REORD_UNIT_71 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_71 ,
										MUX_10_1_IN_1 => UNWINDOWED_71 ,
										MUX_10_1_IN_2 => UNWINDOWED_71 ,
										MUX_10_1_IN_3 => UNWINDOWED_78 ,
										MUX_10_1_IN_4 => UNWINDOWED_78 ,
										MUX_10_1_IN_5 => UNWINDOWED_78 ,
										MUX_10_1_IN_6 => UNWINDOWED_15 ,
										MUX_10_1_IN_7 => UNWINDOWED_142 ,
										MUX_10_1_IN_8 => UNWINDOWED_142 ,
										MUX_10_1_IN_9 => UNWINDOWED_142 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_71
									);
MUX_REORD_UNIT_72 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_72 ,
										MUX_10_1_IN_1 => UNWINDOWED_72 ,
										MUX_10_1_IN_2 => UNWINDOWED_72 ,
										MUX_10_1_IN_3 => UNWINDOWED_65 ,
										MUX_10_1_IN_4 => UNWINDOWED_80 ,
										MUX_10_1_IN_5 => UNWINDOWED_80 ,
										MUX_10_1_IN_6 => UNWINDOWED_17 ,
										MUX_10_1_IN_7 => UNWINDOWED_144 ,
										MUX_10_1_IN_8 => UNWINDOWED_144 ,
										MUX_10_1_IN_9 => UNWINDOWED_144 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_72
									);
MUX_REORD_UNIT_73 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_73 ,
										MUX_10_1_IN_1 => UNWINDOWED_74 ,
										MUX_10_1_IN_2 => UNWINDOWED_74 ,
										MUX_10_1_IN_3 => UNWINDOWED_67 ,
										MUX_10_1_IN_4 => UNWINDOWED_82 ,
										MUX_10_1_IN_5 => UNWINDOWED_82 ,
										MUX_10_1_IN_6 => UNWINDOWED_19 ,
										MUX_10_1_IN_7 => UNWINDOWED_146 ,
										MUX_10_1_IN_8 => UNWINDOWED_146 ,
										MUX_10_1_IN_9 => UNWINDOWED_146 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_73
									);
MUX_REORD_UNIT_74 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_74 ,
										MUX_10_1_IN_1 => UNWINDOWED_73 ,
										MUX_10_1_IN_2 => UNWINDOWED_76 ,
										MUX_10_1_IN_3 => UNWINDOWED_69 ,
										MUX_10_1_IN_4 => UNWINDOWED_84 ,
										MUX_10_1_IN_5 => UNWINDOWED_84 ,
										MUX_10_1_IN_6 => UNWINDOWED_21 ,
										MUX_10_1_IN_7 => UNWINDOWED_148 ,
										MUX_10_1_IN_8 => UNWINDOWED_148 ,
										MUX_10_1_IN_9 => UNWINDOWED_148 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_74
									);
MUX_REORD_UNIT_75 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_75 ,
										MUX_10_1_IN_1 => UNWINDOWED_75 ,
										MUX_10_1_IN_2 => UNWINDOWED_78 ,
										MUX_10_1_IN_3 => UNWINDOWED_71 ,
										MUX_10_1_IN_4 => UNWINDOWED_86 ,
										MUX_10_1_IN_5 => UNWINDOWED_86 ,
										MUX_10_1_IN_6 => UNWINDOWED_23 ,
										MUX_10_1_IN_7 => UNWINDOWED_150 ,
										MUX_10_1_IN_8 => UNWINDOWED_150 ,
										MUX_10_1_IN_9 => UNWINDOWED_150 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_75
									);
MUX_REORD_UNIT_76 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_76 ,
										MUX_10_1_IN_1 => UNWINDOWED_76 ,
										MUX_10_1_IN_2 => UNWINDOWED_73 ,
										MUX_10_1_IN_3 => UNWINDOWED_73 ,
										MUX_10_1_IN_4 => UNWINDOWED_88 ,
										MUX_10_1_IN_5 => UNWINDOWED_88 ,
										MUX_10_1_IN_6 => UNWINDOWED_25 ,
										MUX_10_1_IN_7 => UNWINDOWED_152 ,
										MUX_10_1_IN_8 => UNWINDOWED_152 ,
										MUX_10_1_IN_9 => UNWINDOWED_152 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_76
									);
MUX_REORD_UNIT_77 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_77 ,
										MUX_10_1_IN_1 => UNWINDOWED_78 ,
										MUX_10_1_IN_2 => UNWINDOWED_75 ,
										MUX_10_1_IN_3 => UNWINDOWED_75 ,
										MUX_10_1_IN_4 => UNWINDOWED_90 ,
										MUX_10_1_IN_5 => UNWINDOWED_90 ,
										MUX_10_1_IN_6 => UNWINDOWED_27 ,
										MUX_10_1_IN_7 => UNWINDOWED_154 ,
										MUX_10_1_IN_8 => UNWINDOWED_154 ,
										MUX_10_1_IN_9 => UNWINDOWED_154 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_77
									);
MUX_REORD_UNIT_78 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_78 ,
										MUX_10_1_IN_1 => UNWINDOWED_77 ,
										MUX_10_1_IN_2 => UNWINDOWED_77 ,
										MUX_10_1_IN_3 => UNWINDOWED_77 ,
										MUX_10_1_IN_4 => UNWINDOWED_92 ,
										MUX_10_1_IN_5 => UNWINDOWED_92 ,
										MUX_10_1_IN_6 => UNWINDOWED_29 ,
										MUX_10_1_IN_7 => UNWINDOWED_156 ,
										MUX_10_1_IN_8 => UNWINDOWED_156 ,
										MUX_10_1_IN_9 => UNWINDOWED_156 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_78
									);
MUX_REORD_UNIT_79 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_79 ,
										MUX_10_1_IN_1 => UNWINDOWED_79 ,
										MUX_10_1_IN_2 => UNWINDOWED_79 ,
										MUX_10_1_IN_3 => UNWINDOWED_79 ,
										MUX_10_1_IN_4 => UNWINDOWED_94 ,
										MUX_10_1_IN_5 => UNWINDOWED_94 ,
										MUX_10_1_IN_6 => UNWINDOWED_31 ,
										MUX_10_1_IN_7 => UNWINDOWED_158 ,
										MUX_10_1_IN_8 => UNWINDOWED_158 ,
										MUX_10_1_IN_9 => UNWINDOWED_158 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_79
									);
MUX_REORD_UNIT_80 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_80 ,
										MUX_10_1_IN_1 => UNWINDOWED_80 ,
										MUX_10_1_IN_2 => UNWINDOWED_80 ,
										MUX_10_1_IN_3 => UNWINDOWED_80 ,
										MUX_10_1_IN_4 => UNWINDOWED_65 ,
										MUX_10_1_IN_5 => UNWINDOWED_96 ,
										MUX_10_1_IN_6 => UNWINDOWED_33 ,
										MUX_10_1_IN_7 => UNWINDOWED_160 ,
										MUX_10_1_IN_8 => UNWINDOWED_160 ,
										MUX_10_1_IN_9 => UNWINDOWED_160 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_80
									);
MUX_REORD_UNIT_81 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_81 ,
										MUX_10_1_IN_1 => UNWINDOWED_82 ,
										MUX_10_1_IN_2 => UNWINDOWED_82 ,
										MUX_10_1_IN_3 => UNWINDOWED_82 ,
										MUX_10_1_IN_4 => UNWINDOWED_67 ,
										MUX_10_1_IN_5 => UNWINDOWED_98 ,
										MUX_10_1_IN_6 => UNWINDOWED_35 ,
										MUX_10_1_IN_7 => UNWINDOWED_162 ,
										MUX_10_1_IN_8 => UNWINDOWED_162 ,
										MUX_10_1_IN_9 => UNWINDOWED_162 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_81
									);
MUX_REORD_UNIT_82 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_82 ,
										MUX_10_1_IN_1 => UNWINDOWED_81 ,
										MUX_10_1_IN_2 => UNWINDOWED_84 ,
										MUX_10_1_IN_3 => UNWINDOWED_84 ,
										MUX_10_1_IN_4 => UNWINDOWED_69 ,
										MUX_10_1_IN_5 => UNWINDOWED_100 ,
										MUX_10_1_IN_6 => UNWINDOWED_37 ,
										MUX_10_1_IN_7 => UNWINDOWED_164 ,
										MUX_10_1_IN_8 => UNWINDOWED_164 ,
										MUX_10_1_IN_9 => UNWINDOWED_164 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_82
									);
MUX_REORD_UNIT_83 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_83 ,
										MUX_10_1_IN_1 => UNWINDOWED_83 ,
										MUX_10_1_IN_2 => UNWINDOWED_86 ,
										MUX_10_1_IN_3 => UNWINDOWED_86 ,
										MUX_10_1_IN_4 => UNWINDOWED_71 ,
										MUX_10_1_IN_5 => UNWINDOWED_102 ,
										MUX_10_1_IN_6 => UNWINDOWED_39 ,
										MUX_10_1_IN_7 => UNWINDOWED_166 ,
										MUX_10_1_IN_8 => UNWINDOWED_166 ,
										MUX_10_1_IN_9 => UNWINDOWED_166 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_83
									);
MUX_REORD_UNIT_84 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_84 ,
										MUX_10_1_IN_1 => UNWINDOWED_84 ,
										MUX_10_1_IN_2 => UNWINDOWED_81 ,
										MUX_10_1_IN_3 => UNWINDOWED_88 ,
										MUX_10_1_IN_4 => UNWINDOWED_73 ,
										MUX_10_1_IN_5 => UNWINDOWED_104 ,
										MUX_10_1_IN_6 => UNWINDOWED_41 ,
										MUX_10_1_IN_7 => UNWINDOWED_168 ,
										MUX_10_1_IN_8 => UNWINDOWED_168 ,
										MUX_10_1_IN_9 => UNWINDOWED_168 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_84
									);
MUX_REORD_UNIT_85 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_85 ,
										MUX_10_1_IN_1 => UNWINDOWED_86 ,
										MUX_10_1_IN_2 => UNWINDOWED_83 ,
										MUX_10_1_IN_3 => UNWINDOWED_90 ,
										MUX_10_1_IN_4 => UNWINDOWED_75 ,
										MUX_10_1_IN_5 => UNWINDOWED_106 ,
										MUX_10_1_IN_6 => UNWINDOWED_43 ,
										MUX_10_1_IN_7 => UNWINDOWED_170 ,
										MUX_10_1_IN_8 => UNWINDOWED_170 ,
										MUX_10_1_IN_9 => UNWINDOWED_170 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_85
									);
MUX_REORD_UNIT_86 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_86 ,
										MUX_10_1_IN_1 => UNWINDOWED_85 ,
										MUX_10_1_IN_2 => UNWINDOWED_85 ,
										MUX_10_1_IN_3 => UNWINDOWED_92 ,
										MUX_10_1_IN_4 => UNWINDOWED_77 ,
										MUX_10_1_IN_5 => UNWINDOWED_108 ,
										MUX_10_1_IN_6 => UNWINDOWED_45 ,
										MUX_10_1_IN_7 => UNWINDOWED_172 ,
										MUX_10_1_IN_8 => UNWINDOWED_172 ,
										MUX_10_1_IN_9 => UNWINDOWED_172 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_86
									);
MUX_REORD_UNIT_87 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_87 ,
										MUX_10_1_IN_1 => UNWINDOWED_87 ,
										MUX_10_1_IN_2 => UNWINDOWED_87 ,
										MUX_10_1_IN_3 => UNWINDOWED_94 ,
										MUX_10_1_IN_4 => UNWINDOWED_79 ,
										MUX_10_1_IN_5 => UNWINDOWED_110 ,
										MUX_10_1_IN_6 => UNWINDOWED_47 ,
										MUX_10_1_IN_7 => UNWINDOWED_174 ,
										MUX_10_1_IN_8 => UNWINDOWED_174 ,
										MUX_10_1_IN_9 => UNWINDOWED_174 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_87
									);
MUX_REORD_UNIT_88 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_88 ,
										MUX_10_1_IN_1 => UNWINDOWED_88 ,
										MUX_10_1_IN_2 => UNWINDOWED_88 ,
										MUX_10_1_IN_3 => UNWINDOWED_81 ,
										MUX_10_1_IN_4 => UNWINDOWED_81 ,
										MUX_10_1_IN_5 => UNWINDOWED_112 ,
										MUX_10_1_IN_6 => UNWINDOWED_49 ,
										MUX_10_1_IN_7 => UNWINDOWED_176 ,
										MUX_10_1_IN_8 => UNWINDOWED_176 ,
										MUX_10_1_IN_9 => UNWINDOWED_176 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_88
									);
MUX_REORD_UNIT_89 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_89 ,
										MUX_10_1_IN_1 => UNWINDOWED_90 ,
										MUX_10_1_IN_2 => UNWINDOWED_90 ,
										MUX_10_1_IN_3 => UNWINDOWED_83 ,
										MUX_10_1_IN_4 => UNWINDOWED_83 ,
										MUX_10_1_IN_5 => UNWINDOWED_114 ,
										MUX_10_1_IN_6 => UNWINDOWED_51 ,
										MUX_10_1_IN_7 => UNWINDOWED_178 ,
										MUX_10_1_IN_8 => UNWINDOWED_178 ,
										MUX_10_1_IN_9 => UNWINDOWED_178 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_89
									);
MUX_REORD_UNIT_90 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_90 ,
										MUX_10_1_IN_1 => UNWINDOWED_89 ,
										MUX_10_1_IN_2 => UNWINDOWED_92 ,
										MUX_10_1_IN_3 => UNWINDOWED_85 ,
										MUX_10_1_IN_4 => UNWINDOWED_85 ,
										MUX_10_1_IN_5 => UNWINDOWED_116 ,
										MUX_10_1_IN_6 => UNWINDOWED_53 ,
										MUX_10_1_IN_7 => UNWINDOWED_180 ,
										MUX_10_1_IN_8 => UNWINDOWED_180 ,
										MUX_10_1_IN_9 => UNWINDOWED_180 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_90
									);
MUX_REORD_UNIT_91 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_91 ,
										MUX_10_1_IN_1 => UNWINDOWED_91 ,
										MUX_10_1_IN_2 => UNWINDOWED_94 ,
										MUX_10_1_IN_3 => UNWINDOWED_87 ,
										MUX_10_1_IN_4 => UNWINDOWED_87 ,
										MUX_10_1_IN_5 => UNWINDOWED_118 ,
										MUX_10_1_IN_6 => UNWINDOWED_55 ,
										MUX_10_1_IN_7 => UNWINDOWED_182 ,
										MUX_10_1_IN_8 => UNWINDOWED_182 ,
										MUX_10_1_IN_9 => UNWINDOWED_182 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_91
									);
MUX_REORD_UNIT_92 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_92 ,
										MUX_10_1_IN_1 => UNWINDOWED_92 ,
										MUX_10_1_IN_2 => UNWINDOWED_89 ,
										MUX_10_1_IN_3 => UNWINDOWED_89 ,
										MUX_10_1_IN_4 => UNWINDOWED_89 ,
										MUX_10_1_IN_5 => UNWINDOWED_120 ,
										MUX_10_1_IN_6 => UNWINDOWED_57 ,
										MUX_10_1_IN_7 => UNWINDOWED_184 ,
										MUX_10_1_IN_8 => UNWINDOWED_184 ,
										MUX_10_1_IN_9 => UNWINDOWED_184 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_92
									);
MUX_REORD_UNIT_93 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_93 ,
										MUX_10_1_IN_1 => UNWINDOWED_94 ,
										MUX_10_1_IN_2 => UNWINDOWED_91 ,
										MUX_10_1_IN_3 => UNWINDOWED_91 ,
										MUX_10_1_IN_4 => UNWINDOWED_91 ,
										MUX_10_1_IN_5 => UNWINDOWED_122 ,
										MUX_10_1_IN_6 => UNWINDOWED_59 ,
										MUX_10_1_IN_7 => UNWINDOWED_186 ,
										MUX_10_1_IN_8 => UNWINDOWED_186 ,
										MUX_10_1_IN_9 => UNWINDOWED_186 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_93
									);
MUX_REORD_UNIT_94 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_94 ,
										MUX_10_1_IN_1 => UNWINDOWED_93 ,
										MUX_10_1_IN_2 => UNWINDOWED_93 ,
										MUX_10_1_IN_3 => UNWINDOWED_93 ,
										MUX_10_1_IN_4 => UNWINDOWED_93 ,
										MUX_10_1_IN_5 => UNWINDOWED_124 ,
										MUX_10_1_IN_6 => UNWINDOWED_61 ,
										MUX_10_1_IN_7 => UNWINDOWED_188 ,
										MUX_10_1_IN_8 => UNWINDOWED_188 ,
										MUX_10_1_IN_9 => UNWINDOWED_188 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_94
									);
MUX_REORD_UNIT_95 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_95 ,
										MUX_10_1_IN_1 => UNWINDOWED_95 ,
										MUX_10_1_IN_2 => UNWINDOWED_95 ,
										MUX_10_1_IN_3 => UNWINDOWED_95 ,
										MUX_10_1_IN_4 => UNWINDOWED_95 ,
										MUX_10_1_IN_5 => UNWINDOWED_126 ,
										MUX_10_1_IN_6 => UNWINDOWED_63 ,
										MUX_10_1_IN_7 => UNWINDOWED_190 ,
										MUX_10_1_IN_8 => UNWINDOWED_190 ,
										MUX_10_1_IN_9 => UNWINDOWED_190 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_95
									);
MUX_REORD_UNIT_96 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_96 ,
										MUX_10_1_IN_1 => UNWINDOWED_96 ,
										MUX_10_1_IN_2 => UNWINDOWED_96 ,
										MUX_10_1_IN_3 => UNWINDOWED_96 ,
										MUX_10_1_IN_4 => UNWINDOWED_96 ,
										MUX_10_1_IN_5 => UNWINDOWED_65 ,
										MUX_10_1_IN_6 => UNWINDOWED_65 ,
										MUX_10_1_IN_7 => UNWINDOWED_192 ,
										MUX_10_1_IN_8 => UNWINDOWED_192 ,
										MUX_10_1_IN_9 => UNWINDOWED_192 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_96
									);
MUX_REORD_UNIT_97 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_97 ,
										MUX_10_1_IN_1 => UNWINDOWED_98 ,
										MUX_10_1_IN_2 => UNWINDOWED_98 ,
										MUX_10_1_IN_3 => UNWINDOWED_98 ,
										MUX_10_1_IN_4 => UNWINDOWED_98 ,
										MUX_10_1_IN_5 => UNWINDOWED_67 ,
										MUX_10_1_IN_6 => UNWINDOWED_67 ,
										MUX_10_1_IN_7 => UNWINDOWED_194 ,
										MUX_10_1_IN_8 => UNWINDOWED_194 ,
										MUX_10_1_IN_9 => UNWINDOWED_194 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_97
									);
MUX_REORD_UNIT_98 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_98 ,
										MUX_10_1_IN_1 => UNWINDOWED_97 ,
										MUX_10_1_IN_2 => UNWINDOWED_100 ,
										MUX_10_1_IN_3 => UNWINDOWED_100 ,
										MUX_10_1_IN_4 => UNWINDOWED_100 ,
										MUX_10_1_IN_5 => UNWINDOWED_69 ,
										MUX_10_1_IN_6 => UNWINDOWED_69 ,
										MUX_10_1_IN_7 => UNWINDOWED_196 ,
										MUX_10_1_IN_8 => UNWINDOWED_196 ,
										MUX_10_1_IN_9 => UNWINDOWED_196 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_98
									);
MUX_REORD_UNIT_99 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_99 ,
										MUX_10_1_IN_1 => UNWINDOWED_99 ,
										MUX_10_1_IN_2 => UNWINDOWED_102 ,
										MUX_10_1_IN_3 => UNWINDOWED_102 ,
										MUX_10_1_IN_4 => UNWINDOWED_102 ,
										MUX_10_1_IN_5 => UNWINDOWED_71 ,
										MUX_10_1_IN_6 => UNWINDOWED_71 ,
										MUX_10_1_IN_7 => UNWINDOWED_198 ,
										MUX_10_1_IN_8 => UNWINDOWED_198 ,
										MUX_10_1_IN_9 => UNWINDOWED_198 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_99
									);
MUX_REORD_UNIT_100 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_100 ,
										MUX_10_1_IN_1 => UNWINDOWED_100 ,
										MUX_10_1_IN_2 => UNWINDOWED_97 ,
										MUX_10_1_IN_3 => UNWINDOWED_104 ,
										MUX_10_1_IN_4 => UNWINDOWED_104 ,
										MUX_10_1_IN_5 => UNWINDOWED_73 ,
										MUX_10_1_IN_6 => UNWINDOWED_73 ,
										MUX_10_1_IN_7 => UNWINDOWED_200 ,
										MUX_10_1_IN_8 => UNWINDOWED_200 ,
										MUX_10_1_IN_9 => UNWINDOWED_200 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_100
									);
MUX_REORD_UNIT_101 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_101 ,
										MUX_10_1_IN_1 => UNWINDOWED_102 ,
										MUX_10_1_IN_2 => UNWINDOWED_99 ,
										MUX_10_1_IN_3 => UNWINDOWED_106 ,
										MUX_10_1_IN_4 => UNWINDOWED_106 ,
										MUX_10_1_IN_5 => UNWINDOWED_75 ,
										MUX_10_1_IN_6 => UNWINDOWED_75 ,
										MUX_10_1_IN_7 => UNWINDOWED_202 ,
										MUX_10_1_IN_8 => UNWINDOWED_202 ,
										MUX_10_1_IN_9 => UNWINDOWED_202 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_101
									);
MUX_REORD_UNIT_102 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_102 ,
										MUX_10_1_IN_1 => UNWINDOWED_101 ,
										MUX_10_1_IN_2 => UNWINDOWED_101 ,
										MUX_10_1_IN_3 => UNWINDOWED_108 ,
										MUX_10_1_IN_4 => UNWINDOWED_108 ,
										MUX_10_1_IN_5 => UNWINDOWED_77 ,
										MUX_10_1_IN_6 => UNWINDOWED_77 ,
										MUX_10_1_IN_7 => UNWINDOWED_204 ,
										MUX_10_1_IN_8 => UNWINDOWED_204 ,
										MUX_10_1_IN_9 => UNWINDOWED_204 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_102
									);
MUX_REORD_UNIT_103 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_103 ,
										MUX_10_1_IN_1 => UNWINDOWED_103 ,
										MUX_10_1_IN_2 => UNWINDOWED_103 ,
										MUX_10_1_IN_3 => UNWINDOWED_110 ,
										MUX_10_1_IN_4 => UNWINDOWED_110 ,
										MUX_10_1_IN_5 => UNWINDOWED_79 ,
										MUX_10_1_IN_6 => UNWINDOWED_79 ,
										MUX_10_1_IN_7 => UNWINDOWED_206 ,
										MUX_10_1_IN_8 => UNWINDOWED_206 ,
										MUX_10_1_IN_9 => UNWINDOWED_206 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_103
									);
MUX_REORD_UNIT_104 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_104 ,
										MUX_10_1_IN_1 => UNWINDOWED_104 ,
										MUX_10_1_IN_2 => UNWINDOWED_104 ,
										MUX_10_1_IN_3 => UNWINDOWED_97 ,
										MUX_10_1_IN_4 => UNWINDOWED_112 ,
										MUX_10_1_IN_5 => UNWINDOWED_81 ,
										MUX_10_1_IN_6 => UNWINDOWED_81 ,
										MUX_10_1_IN_7 => UNWINDOWED_208 ,
										MUX_10_1_IN_8 => UNWINDOWED_208 ,
										MUX_10_1_IN_9 => UNWINDOWED_208 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_104
									);
MUX_REORD_UNIT_105 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_105 ,
										MUX_10_1_IN_1 => UNWINDOWED_106 ,
										MUX_10_1_IN_2 => UNWINDOWED_106 ,
										MUX_10_1_IN_3 => UNWINDOWED_99 ,
										MUX_10_1_IN_4 => UNWINDOWED_114 ,
										MUX_10_1_IN_5 => UNWINDOWED_83 ,
										MUX_10_1_IN_6 => UNWINDOWED_83 ,
										MUX_10_1_IN_7 => UNWINDOWED_210 ,
										MUX_10_1_IN_8 => UNWINDOWED_210 ,
										MUX_10_1_IN_9 => UNWINDOWED_210 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_105
									);
MUX_REORD_UNIT_106 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_106 ,
										MUX_10_1_IN_1 => UNWINDOWED_105 ,
										MUX_10_1_IN_2 => UNWINDOWED_108 ,
										MUX_10_1_IN_3 => UNWINDOWED_101 ,
										MUX_10_1_IN_4 => UNWINDOWED_116 ,
										MUX_10_1_IN_5 => UNWINDOWED_85 ,
										MUX_10_1_IN_6 => UNWINDOWED_85 ,
										MUX_10_1_IN_7 => UNWINDOWED_212 ,
										MUX_10_1_IN_8 => UNWINDOWED_212 ,
										MUX_10_1_IN_9 => UNWINDOWED_212 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_106
									);
MUX_REORD_UNIT_107 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_107 ,
										MUX_10_1_IN_1 => UNWINDOWED_107 ,
										MUX_10_1_IN_2 => UNWINDOWED_110 ,
										MUX_10_1_IN_3 => UNWINDOWED_103 ,
										MUX_10_1_IN_4 => UNWINDOWED_118 ,
										MUX_10_1_IN_5 => UNWINDOWED_87 ,
										MUX_10_1_IN_6 => UNWINDOWED_87 ,
										MUX_10_1_IN_7 => UNWINDOWED_214 ,
										MUX_10_1_IN_8 => UNWINDOWED_214 ,
										MUX_10_1_IN_9 => UNWINDOWED_214 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_107
									);
MUX_REORD_UNIT_108 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_108 ,
										MUX_10_1_IN_1 => UNWINDOWED_108 ,
										MUX_10_1_IN_2 => UNWINDOWED_105 ,
										MUX_10_1_IN_3 => UNWINDOWED_105 ,
										MUX_10_1_IN_4 => UNWINDOWED_120 ,
										MUX_10_1_IN_5 => UNWINDOWED_89 ,
										MUX_10_1_IN_6 => UNWINDOWED_89 ,
										MUX_10_1_IN_7 => UNWINDOWED_216 ,
										MUX_10_1_IN_8 => UNWINDOWED_216 ,
										MUX_10_1_IN_9 => UNWINDOWED_216 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_108
									);
MUX_REORD_UNIT_109 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_109 ,
										MUX_10_1_IN_1 => UNWINDOWED_110 ,
										MUX_10_1_IN_2 => UNWINDOWED_107 ,
										MUX_10_1_IN_3 => UNWINDOWED_107 ,
										MUX_10_1_IN_4 => UNWINDOWED_122 ,
										MUX_10_1_IN_5 => UNWINDOWED_91 ,
										MUX_10_1_IN_6 => UNWINDOWED_91 ,
										MUX_10_1_IN_7 => UNWINDOWED_218 ,
										MUX_10_1_IN_8 => UNWINDOWED_218 ,
										MUX_10_1_IN_9 => UNWINDOWED_218 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_109
									);
MUX_REORD_UNIT_110 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_110 ,
										MUX_10_1_IN_1 => UNWINDOWED_109 ,
										MUX_10_1_IN_2 => UNWINDOWED_109 ,
										MUX_10_1_IN_3 => UNWINDOWED_109 ,
										MUX_10_1_IN_4 => UNWINDOWED_124 ,
										MUX_10_1_IN_5 => UNWINDOWED_93 ,
										MUX_10_1_IN_6 => UNWINDOWED_93 ,
										MUX_10_1_IN_7 => UNWINDOWED_220 ,
										MUX_10_1_IN_8 => UNWINDOWED_220 ,
										MUX_10_1_IN_9 => UNWINDOWED_220 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_110
									);
MUX_REORD_UNIT_111 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_111 ,
										MUX_10_1_IN_1 => UNWINDOWED_111 ,
										MUX_10_1_IN_2 => UNWINDOWED_111 ,
										MUX_10_1_IN_3 => UNWINDOWED_111 ,
										MUX_10_1_IN_4 => UNWINDOWED_126 ,
										MUX_10_1_IN_5 => UNWINDOWED_95 ,
										MUX_10_1_IN_6 => UNWINDOWED_95 ,
										MUX_10_1_IN_7 => UNWINDOWED_222 ,
										MUX_10_1_IN_8 => UNWINDOWED_222 ,
										MUX_10_1_IN_9 => UNWINDOWED_222 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_111
									);
MUX_REORD_UNIT_112 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_112 ,
										MUX_10_1_IN_1 => UNWINDOWED_112 ,
										MUX_10_1_IN_2 => UNWINDOWED_112 ,
										MUX_10_1_IN_3 => UNWINDOWED_112 ,
										MUX_10_1_IN_4 => UNWINDOWED_97 ,
										MUX_10_1_IN_5 => UNWINDOWED_97 ,
										MUX_10_1_IN_6 => UNWINDOWED_97 ,
										MUX_10_1_IN_7 => UNWINDOWED_224 ,
										MUX_10_1_IN_8 => UNWINDOWED_224 ,
										MUX_10_1_IN_9 => UNWINDOWED_224 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_112
									);
MUX_REORD_UNIT_113 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_113 ,
										MUX_10_1_IN_1 => UNWINDOWED_114 ,
										MUX_10_1_IN_2 => UNWINDOWED_114 ,
										MUX_10_1_IN_3 => UNWINDOWED_114 ,
										MUX_10_1_IN_4 => UNWINDOWED_99 ,
										MUX_10_1_IN_5 => UNWINDOWED_99 ,
										MUX_10_1_IN_6 => UNWINDOWED_99 ,
										MUX_10_1_IN_7 => UNWINDOWED_226 ,
										MUX_10_1_IN_8 => UNWINDOWED_226 ,
										MUX_10_1_IN_9 => UNWINDOWED_226 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_113
									);
MUX_REORD_UNIT_114 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_114 ,
										MUX_10_1_IN_1 => UNWINDOWED_113 ,
										MUX_10_1_IN_2 => UNWINDOWED_116 ,
										MUX_10_1_IN_3 => UNWINDOWED_116 ,
										MUX_10_1_IN_4 => UNWINDOWED_101 ,
										MUX_10_1_IN_5 => UNWINDOWED_101 ,
										MUX_10_1_IN_6 => UNWINDOWED_101 ,
										MUX_10_1_IN_7 => UNWINDOWED_228 ,
										MUX_10_1_IN_8 => UNWINDOWED_228 ,
										MUX_10_1_IN_9 => UNWINDOWED_228 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_114
									);
MUX_REORD_UNIT_115 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_115 ,
										MUX_10_1_IN_1 => UNWINDOWED_115 ,
										MUX_10_1_IN_2 => UNWINDOWED_118 ,
										MUX_10_1_IN_3 => UNWINDOWED_118 ,
										MUX_10_1_IN_4 => UNWINDOWED_103 ,
										MUX_10_1_IN_5 => UNWINDOWED_103 ,
										MUX_10_1_IN_6 => UNWINDOWED_103 ,
										MUX_10_1_IN_7 => UNWINDOWED_230 ,
										MUX_10_1_IN_8 => UNWINDOWED_230 ,
										MUX_10_1_IN_9 => UNWINDOWED_230 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_115
									);
MUX_REORD_UNIT_116 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_116 ,
										MUX_10_1_IN_1 => UNWINDOWED_116 ,
										MUX_10_1_IN_2 => UNWINDOWED_113 ,
										MUX_10_1_IN_3 => UNWINDOWED_120 ,
										MUX_10_1_IN_4 => UNWINDOWED_105 ,
										MUX_10_1_IN_5 => UNWINDOWED_105 ,
										MUX_10_1_IN_6 => UNWINDOWED_105 ,
										MUX_10_1_IN_7 => UNWINDOWED_232 ,
										MUX_10_1_IN_8 => UNWINDOWED_232 ,
										MUX_10_1_IN_9 => UNWINDOWED_232 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_116
									);
MUX_REORD_UNIT_117 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_117 ,
										MUX_10_1_IN_1 => UNWINDOWED_118 ,
										MUX_10_1_IN_2 => UNWINDOWED_115 ,
										MUX_10_1_IN_3 => UNWINDOWED_122 ,
										MUX_10_1_IN_4 => UNWINDOWED_107 ,
										MUX_10_1_IN_5 => UNWINDOWED_107 ,
										MUX_10_1_IN_6 => UNWINDOWED_107 ,
										MUX_10_1_IN_7 => UNWINDOWED_234 ,
										MUX_10_1_IN_8 => UNWINDOWED_234 ,
										MUX_10_1_IN_9 => UNWINDOWED_234 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_117
									);
MUX_REORD_UNIT_118 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_118 ,
										MUX_10_1_IN_1 => UNWINDOWED_117 ,
										MUX_10_1_IN_2 => UNWINDOWED_117 ,
										MUX_10_1_IN_3 => UNWINDOWED_124 ,
										MUX_10_1_IN_4 => UNWINDOWED_109 ,
										MUX_10_1_IN_5 => UNWINDOWED_109 ,
										MUX_10_1_IN_6 => UNWINDOWED_109 ,
										MUX_10_1_IN_7 => UNWINDOWED_236 ,
										MUX_10_1_IN_8 => UNWINDOWED_236 ,
										MUX_10_1_IN_9 => UNWINDOWED_236 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_118
									);
MUX_REORD_UNIT_119 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_119 ,
										MUX_10_1_IN_1 => UNWINDOWED_119 ,
										MUX_10_1_IN_2 => UNWINDOWED_119 ,
										MUX_10_1_IN_3 => UNWINDOWED_126 ,
										MUX_10_1_IN_4 => UNWINDOWED_111 ,
										MUX_10_1_IN_5 => UNWINDOWED_111 ,
										MUX_10_1_IN_6 => UNWINDOWED_111 ,
										MUX_10_1_IN_7 => UNWINDOWED_238 ,
										MUX_10_1_IN_8 => UNWINDOWED_238 ,
										MUX_10_1_IN_9 => UNWINDOWED_238 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_119
									);
MUX_REORD_UNIT_120 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_120 ,
										MUX_10_1_IN_1 => UNWINDOWED_120 ,
										MUX_10_1_IN_2 => UNWINDOWED_120 ,
										MUX_10_1_IN_3 => UNWINDOWED_113 ,
										MUX_10_1_IN_4 => UNWINDOWED_113 ,
										MUX_10_1_IN_5 => UNWINDOWED_113 ,
										MUX_10_1_IN_6 => UNWINDOWED_113 ,
										MUX_10_1_IN_7 => UNWINDOWED_240 ,
										MUX_10_1_IN_8 => UNWINDOWED_240 ,
										MUX_10_1_IN_9 => UNWINDOWED_240 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_120
									);
MUX_REORD_UNIT_121 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_121 ,
										MUX_10_1_IN_1 => UNWINDOWED_122 ,
										MUX_10_1_IN_2 => UNWINDOWED_122 ,
										MUX_10_1_IN_3 => UNWINDOWED_115 ,
										MUX_10_1_IN_4 => UNWINDOWED_115 ,
										MUX_10_1_IN_5 => UNWINDOWED_115 ,
										MUX_10_1_IN_6 => UNWINDOWED_115 ,
										MUX_10_1_IN_7 => UNWINDOWED_242 ,
										MUX_10_1_IN_8 => UNWINDOWED_242 ,
										MUX_10_1_IN_9 => UNWINDOWED_242 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_121
									);
MUX_REORD_UNIT_122 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_122 ,
										MUX_10_1_IN_1 => UNWINDOWED_121 ,
										MUX_10_1_IN_2 => UNWINDOWED_124 ,
										MUX_10_1_IN_3 => UNWINDOWED_117 ,
										MUX_10_1_IN_4 => UNWINDOWED_117 ,
										MUX_10_1_IN_5 => UNWINDOWED_117 ,
										MUX_10_1_IN_6 => UNWINDOWED_117 ,
										MUX_10_1_IN_7 => UNWINDOWED_244 ,
										MUX_10_1_IN_8 => UNWINDOWED_244 ,
										MUX_10_1_IN_9 => UNWINDOWED_244 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_122
									);
MUX_REORD_UNIT_123 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_123 ,
										MUX_10_1_IN_1 => UNWINDOWED_123 ,
										MUX_10_1_IN_2 => UNWINDOWED_126 ,
										MUX_10_1_IN_3 => UNWINDOWED_119 ,
										MUX_10_1_IN_4 => UNWINDOWED_119 ,
										MUX_10_1_IN_5 => UNWINDOWED_119 ,
										MUX_10_1_IN_6 => UNWINDOWED_119 ,
										MUX_10_1_IN_7 => UNWINDOWED_246 ,
										MUX_10_1_IN_8 => UNWINDOWED_246 ,
										MUX_10_1_IN_9 => UNWINDOWED_246 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_123
									);
MUX_REORD_UNIT_124 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_124 ,
										MUX_10_1_IN_1 => UNWINDOWED_124 ,
										MUX_10_1_IN_2 => UNWINDOWED_121 ,
										MUX_10_1_IN_3 => UNWINDOWED_121 ,
										MUX_10_1_IN_4 => UNWINDOWED_121 ,
										MUX_10_1_IN_5 => UNWINDOWED_121 ,
										MUX_10_1_IN_6 => UNWINDOWED_121 ,
										MUX_10_1_IN_7 => UNWINDOWED_248 ,
										MUX_10_1_IN_8 => UNWINDOWED_248 ,
										MUX_10_1_IN_9 => UNWINDOWED_248 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_124
									);
MUX_REORD_UNIT_125 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_125 ,
										MUX_10_1_IN_1 => UNWINDOWED_126 ,
										MUX_10_1_IN_2 => UNWINDOWED_123 ,
										MUX_10_1_IN_3 => UNWINDOWED_123 ,
										MUX_10_1_IN_4 => UNWINDOWED_123 ,
										MUX_10_1_IN_5 => UNWINDOWED_123 ,
										MUX_10_1_IN_6 => UNWINDOWED_123 ,
										MUX_10_1_IN_7 => UNWINDOWED_250 ,
										MUX_10_1_IN_8 => UNWINDOWED_250 ,
										MUX_10_1_IN_9 => UNWINDOWED_250 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_125
									);
MUX_REORD_UNIT_126 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_126 ,
										MUX_10_1_IN_1 => UNWINDOWED_125 ,
										MUX_10_1_IN_2 => UNWINDOWED_125 ,
										MUX_10_1_IN_3 => UNWINDOWED_125 ,
										MUX_10_1_IN_4 => UNWINDOWED_125 ,
										MUX_10_1_IN_5 => UNWINDOWED_125 ,
										MUX_10_1_IN_6 => UNWINDOWED_125 ,
										MUX_10_1_IN_7 => UNWINDOWED_252 ,
										MUX_10_1_IN_8 => UNWINDOWED_252 ,
										MUX_10_1_IN_9 => UNWINDOWED_252 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_126
									);
MUX_REORD_UNIT_127 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_127 ,
										MUX_10_1_IN_1 => UNWINDOWED_127 ,
										MUX_10_1_IN_2 => UNWINDOWED_127 ,
										MUX_10_1_IN_3 => UNWINDOWED_127 ,
										MUX_10_1_IN_4 => UNWINDOWED_127 ,
										MUX_10_1_IN_5 => UNWINDOWED_127 ,
										MUX_10_1_IN_6 => UNWINDOWED_127 ,
										MUX_10_1_IN_7 => UNWINDOWED_254 ,
										MUX_10_1_IN_8 => UNWINDOWED_254 ,
										MUX_10_1_IN_9 => UNWINDOWED_254 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_127
									);
MUX_REORD_UNIT_128 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_128 ,
										MUX_10_1_IN_1 => UNWINDOWED_128 ,
										MUX_10_1_IN_2 => UNWINDOWED_128 ,
										MUX_10_1_IN_3 => UNWINDOWED_128 ,
										MUX_10_1_IN_4 => UNWINDOWED_128 ,
										MUX_10_1_IN_5 => UNWINDOWED_128 ,
										MUX_10_1_IN_6 => UNWINDOWED_128 ,
										MUX_10_1_IN_7 => UNWINDOWED_1 ,
										MUX_10_1_IN_8 => UNWINDOWED_256 ,
										MUX_10_1_IN_9 => UNWINDOWED_256 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_128
									);
MUX_REORD_UNIT_129 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_129 ,
										MUX_10_1_IN_1 => UNWINDOWED_130 ,
										MUX_10_1_IN_2 => UNWINDOWED_130 ,
										MUX_10_1_IN_3 => UNWINDOWED_130 ,
										MUX_10_1_IN_4 => UNWINDOWED_130 ,
										MUX_10_1_IN_5 => UNWINDOWED_130 ,
										MUX_10_1_IN_6 => UNWINDOWED_130 ,
										MUX_10_1_IN_7 => UNWINDOWED_3 ,
										MUX_10_1_IN_8 => UNWINDOWED_258 ,
										MUX_10_1_IN_9 => UNWINDOWED_258 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_129
									);
MUX_REORD_UNIT_130 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_130 ,
										MUX_10_1_IN_1 => UNWINDOWED_129 ,
										MUX_10_1_IN_2 => UNWINDOWED_132 ,
										MUX_10_1_IN_3 => UNWINDOWED_132 ,
										MUX_10_1_IN_4 => UNWINDOWED_132 ,
										MUX_10_1_IN_5 => UNWINDOWED_132 ,
										MUX_10_1_IN_6 => UNWINDOWED_132 ,
										MUX_10_1_IN_7 => UNWINDOWED_5 ,
										MUX_10_1_IN_8 => UNWINDOWED_260 ,
										MUX_10_1_IN_9 => UNWINDOWED_260 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_130
									);
MUX_REORD_UNIT_131 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_131 ,
										MUX_10_1_IN_1 => UNWINDOWED_131 ,
										MUX_10_1_IN_2 => UNWINDOWED_134 ,
										MUX_10_1_IN_3 => UNWINDOWED_134 ,
										MUX_10_1_IN_4 => UNWINDOWED_134 ,
										MUX_10_1_IN_5 => UNWINDOWED_134 ,
										MUX_10_1_IN_6 => UNWINDOWED_134 ,
										MUX_10_1_IN_7 => UNWINDOWED_7 ,
										MUX_10_1_IN_8 => UNWINDOWED_262 ,
										MUX_10_1_IN_9 => UNWINDOWED_262 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_131
									);
MUX_REORD_UNIT_132 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_132 ,
										MUX_10_1_IN_1 => UNWINDOWED_132 ,
										MUX_10_1_IN_2 => UNWINDOWED_129 ,
										MUX_10_1_IN_3 => UNWINDOWED_136 ,
										MUX_10_1_IN_4 => UNWINDOWED_136 ,
										MUX_10_1_IN_5 => UNWINDOWED_136 ,
										MUX_10_1_IN_6 => UNWINDOWED_136 ,
										MUX_10_1_IN_7 => UNWINDOWED_9 ,
										MUX_10_1_IN_8 => UNWINDOWED_264 ,
										MUX_10_1_IN_9 => UNWINDOWED_264 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_132
									);
MUX_REORD_UNIT_133 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_133 ,
										MUX_10_1_IN_1 => UNWINDOWED_134 ,
										MUX_10_1_IN_2 => UNWINDOWED_131 ,
										MUX_10_1_IN_3 => UNWINDOWED_138 ,
										MUX_10_1_IN_4 => UNWINDOWED_138 ,
										MUX_10_1_IN_5 => UNWINDOWED_138 ,
										MUX_10_1_IN_6 => UNWINDOWED_138 ,
										MUX_10_1_IN_7 => UNWINDOWED_11 ,
										MUX_10_1_IN_8 => UNWINDOWED_266 ,
										MUX_10_1_IN_9 => UNWINDOWED_266 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_133
									);
MUX_REORD_UNIT_134 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_134 ,
										MUX_10_1_IN_1 => UNWINDOWED_133 ,
										MUX_10_1_IN_2 => UNWINDOWED_133 ,
										MUX_10_1_IN_3 => UNWINDOWED_140 ,
										MUX_10_1_IN_4 => UNWINDOWED_140 ,
										MUX_10_1_IN_5 => UNWINDOWED_140 ,
										MUX_10_1_IN_6 => UNWINDOWED_140 ,
										MUX_10_1_IN_7 => UNWINDOWED_13 ,
										MUX_10_1_IN_8 => UNWINDOWED_268 ,
										MUX_10_1_IN_9 => UNWINDOWED_268 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_134
									);
MUX_REORD_UNIT_135 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_135 ,
										MUX_10_1_IN_1 => UNWINDOWED_135 ,
										MUX_10_1_IN_2 => UNWINDOWED_135 ,
										MUX_10_1_IN_3 => UNWINDOWED_142 ,
										MUX_10_1_IN_4 => UNWINDOWED_142 ,
										MUX_10_1_IN_5 => UNWINDOWED_142 ,
										MUX_10_1_IN_6 => UNWINDOWED_142 ,
										MUX_10_1_IN_7 => UNWINDOWED_15 ,
										MUX_10_1_IN_8 => UNWINDOWED_270 ,
										MUX_10_1_IN_9 => UNWINDOWED_270 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_135
									);
MUX_REORD_UNIT_136 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_136 ,
										MUX_10_1_IN_1 => UNWINDOWED_136 ,
										MUX_10_1_IN_2 => UNWINDOWED_136 ,
										MUX_10_1_IN_3 => UNWINDOWED_129 ,
										MUX_10_1_IN_4 => UNWINDOWED_144 ,
										MUX_10_1_IN_5 => UNWINDOWED_144 ,
										MUX_10_1_IN_6 => UNWINDOWED_144 ,
										MUX_10_1_IN_7 => UNWINDOWED_17 ,
										MUX_10_1_IN_8 => UNWINDOWED_272 ,
										MUX_10_1_IN_9 => UNWINDOWED_272 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_136
									);
MUX_REORD_UNIT_137 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_137 ,
										MUX_10_1_IN_1 => UNWINDOWED_138 ,
										MUX_10_1_IN_2 => UNWINDOWED_138 ,
										MUX_10_1_IN_3 => UNWINDOWED_131 ,
										MUX_10_1_IN_4 => UNWINDOWED_146 ,
										MUX_10_1_IN_5 => UNWINDOWED_146 ,
										MUX_10_1_IN_6 => UNWINDOWED_146 ,
										MUX_10_1_IN_7 => UNWINDOWED_19 ,
										MUX_10_1_IN_8 => UNWINDOWED_274 ,
										MUX_10_1_IN_9 => UNWINDOWED_274 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_137
									);
MUX_REORD_UNIT_138 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_138 ,
										MUX_10_1_IN_1 => UNWINDOWED_137 ,
										MUX_10_1_IN_2 => UNWINDOWED_140 ,
										MUX_10_1_IN_3 => UNWINDOWED_133 ,
										MUX_10_1_IN_4 => UNWINDOWED_148 ,
										MUX_10_1_IN_5 => UNWINDOWED_148 ,
										MUX_10_1_IN_6 => UNWINDOWED_148 ,
										MUX_10_1_IN_7 => UNWINDOWED_21 ,
										MUX_10_1_IN_8 => UNWINDOWED_276 ,
										MUX_10_1_IN_9 => UNWINDOWED_276 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_138
									);
MUX_REORD_UNIT_139 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_139 ,
										MUX_10_1_IN_1 => UNWINDOWED_139 ,
										MUX_10_1_IN_2 => UNWINDOWED_142 ,
										MUX_10_1_IN_3 => UNWINDOWED_135 ,
										MUX_10_1_IN_4 => UNWINDOWED_150 ,
										MUX_10_1_IN_5 => UNWINDOWED_150 ,
										MUX_10_1_IN_6 => UNWINDOWED_150 ,
										MUX_10_1_IN_7 => UNWINDOWED_23 ,
										MUX_10_1_IN_8 => UNWINDOWED_278 ,
										MUX_10_1_IN_9 => UNWINDOWED_278 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_139
									);
MUX_REORD_UNIT_140 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_140 ,
										MUX_10_1_IN_1 => UNWINDOWED_140 ,
										MUX_10_1_IN_2 => UNWINDOWED_137 ,
										MUX_10_1_IN_3 => UNWINDOWED_137 ,
										MUX_10_1_IN_4 => UNWINDOWED_152 ,
										MUX_10_1_IN_5 => UNWINDOWED_152 ,
										MUX_10_1_IN_6 => UNWINDOWED_152 ,
										MUX_10_1_IN_7 => UNWINDOWED_25 ,
										MUX_10_1_IN_8 => UNWINDOWED_280 ,
										MUX_10_1_IN_9 => UNWINDOWED_280 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_140
									);
MUX_REORD_UNIT_141 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_141 ,
										MUX_10_1_IN_1 => UNWINDOWED_142 ,
										MUX_10_1_IN_2 => UNWINDOWED_139 ,
										MUX_10_1_IN_3 => UNWINDOWED_139 ,
										MUX_10_1_IN_4 => UNWINDOWED_154 ,
										MUX_10_1_IN_5 => UNWINDOWED_154 ,
										MUX_10_1_IN_6 => UNWINDOWED_154 ,
										MUX_10_1_IN_7 => UNWINDOWED_27 ,
										MUX_10_1_IN_8 => UNWINDOWED_282 ,
										MUX_10_1_IN_9 => UNWINDOWED_282 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_141
									);
MUX_REORD_UNIT_142 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_142 ,
										MUX_10_1_IN_1 => UNWINDOWED_141 ,
										MUX_10_1_IN_2 => UNWINDOWED_141 ,
										MUX_10_1_IN_3 => UNWINDOWED_141 ,
										MUX_10_1_IN_4 => UNWINDOWED_156 ,
										MUX_10_1_IN_5 => UNWINDOWED_156 ,
										MUX_10_1_IN_6 => UNWINDOWED_156 ,
										MUX_10_1_IN_7 => UNWINDOWED_29 ,
										MUX_10_1_IN_8 => UNWINDOWED_284 ,
										MUX_10_1_IN_9 => UNWINDOWED_284 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_142
									);
MUX_REORD_UNIT_143 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_143 ,
										MUX_10_1_IN_1 => UNWINDOWED_143 ,
										MUX_10_1_IN_2 => UNWINDOWED_143 ,
										MUX_10_1_IN_3 => UNWINDOWED_143 ,
										MUX_10_1_IN_4 => UNWINDOWED_158 ,
										MUX_10_1_IN_5 => UNWINDOWED_158 ,
										MUX_10_1_IN_6 => UNWINDOWED_158 ,
										MUX_10_1_IN_7 => UNWINDOWED_31 ,
										MUX_10_1_IN_8 => UNWINDOWED_286 ,
										MUX_10_1_IN_9 => UNWINDOWED_286 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_143
									);
MUX_REORD_UNIT_144 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_144 ,
										MUX_10_1_IN_1 => UNWINDOWED_144 ,
										MUX_10_1_IN_2 => UNWINDOWED_144 ,
										MUX_10_1_IN_3 => UNWINDOWED_144 ,
										MUX_10_1_IN_4 => UNWINDOWED_129 ,
										MUX_10_1_IN_5 => UNWINDOWED_160 ,
										MUX_10_1_IN_6 => UNWINDOWED_160 ,
										MUX_10_1_IN_7 => UNWINDOWED_33 ,
										MUX_10_1_IN_8 => UNWINDOWED_288 ,
										MUX_10_1_IN_9 => UNWINDOWED_288 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_144
									);
MUX_REORD_UNIT_145 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_145 ,
										MUX_10_1_IN_1 => UNWINDOWED_146 ,
										MUX_10_1_IN_2 => UNWINDOWED_146 ,
										MUX_10_1_IN_3 => UNWINDOWED_146 ,
										MUX_10_1_IN_4 => UNWINDOWED_131 ,
										MUX_10_1_IN_5 => UNWINDOWED_162 ,
										MUX_10_1_IN_6 => UNWINDOWED_162 ,
										MUX_10_1_IN_7 => UNWINDOWED_35 ,
										MUX_10_1_IN_8 => UNWINDOWED_290 ,
										MUX_10_1_IN_9 => UNWINDOWED_290 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_145
									);
MUX_REORD_UNIT_146 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_146 ,
										MUX_10_1_IN_1 => UNWINDOWED_145 ,
										MUX_10_1_IN_2 => UNWINDOWED_148 ,
										MUX_10_1_IN_3 => UNWINDOWED_148 ,
										MUX_10_1_IN_4 => UNWINDOWED_133 ,
										MUX_10_1_IN_5 => UNWINDOWED_164 ,
										MUX_10_1_IN_6 => UNWINDOWED_164 ,
										MUX_10_1_IN_7 => UNWINDOWED_37 ,
										MUX_10_1_IN_8 => UNWINDOWED_292 ,
										MUX_10_1_IN_9 => UNWINDOWED_292 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_146
									);
MUX_REORD_UNIT_147 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_147 ,
										MUX_10_1_IN_1 => UNWINDOWED_147 ,
										MUX_10_1_IN_2 => UNWINDOWED_150 ,
										MUX_10_1_IN_3 => UNWINDOWED_150 ,
										MUX_10_1_IN_4 => UNWINDOWED_135 ,
										MUX_10_1_IN_5 => UNWINDOWED_166 ,
										MUX_10_1_IN_6 => UNWINDOWED_166 ,
										MUX_10_1_IN_7 => UNWINDOWED_39 ,
										MUX_10_1_IN_8 => UNWINDOWED_294 ,
										MUX_10_1_IN_9 => UNWINDOWED_294 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_147
									);
MUX_REORD_UNIT_148 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_148 ,
										MUX_10_1_IN_1 => UNWINDOWED_148 ,
										MUX_10_1_IN_2 => UNWINDOWED_145 ,
										MUX_10_1_IN_3 => UNWINDOWED_152 ,
										MUX_10_1_IN_4 => UNWINDOWED_137 ,
										MUX_10_1_IN_5 => UNWINDOWED_168 ,
										MUX_10_1_IN_6 => UNWINDOWED_168 ,
										MUX_10_1_IN_7 => UNWINDOWED_41 ,
										MUX_10_1_IN_8 => UNWINDOWED_296 ,
										MUX_10_1_IN_9 => UNWINDOWED_296 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_148
									);
MUX_REORD_UNIT_149 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_149 ,
										MUX_10_1_IN_1 => UNWINDOWED_150 ,
										MUX_10_1_IN_2 => UNWINDOWED_147 ,
										MUX_10_1_IN_3 => UNWINDOWED_154 ,
										MUX_10_1_IN_4 => UNWINDOWED_139 ,
										MUX_10_1_IN_5 => UNWINDOWED_170 ,
										MUX_10_1_IN_6 => UNWINDOWED_170 ,
										MUX_10_1_IN_7 => UNWINDOWED_43 ,
										MUX_10_1_IN_8 => UNWINDOWED_298 ,
										MUX_10_1_IN_9 => UNWINDOWED_298 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_149
									);
MUX_REORD_UNIT_150 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_150 ,
										MUX_10_1_IN_1 => UNWINDOWED_149 ,
										MUX_10_1_IN_2 => UNWINDOWED_149 ,
										MUX_10_1_IN_3 => UNWINDOWED_156 ,
										MUX_10_1_IN_4 => UNWINDOWED_141 ,
										MUX_10_1_IN_5 => UNWINDOWED_172 ,
										MUX_10_1_IN_6 => UNWINDOWED_172 ,
										MUX_10_1_IN_7 => UNWINDOWED_45 ,
										MUX_10_1_IN_8 => UNWINDOWED_300 ,
										MUX_10_1_IN_9 => UNWINDOWED_300 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_150
									);
MUX_REORD_UNIT_151 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_151 ,
										MUX_10_1_IN_1 => UNWINDOWED_151 ,
										MUX_10_1_IN_2 => UNWINDOWED_151 ,
										MUX_10_1_IN_3 => UNWINDOWED_158 ,
										MUX_10_1_IN_4 => UNWINDOWED_143 ,
										MUX_10_1_IN_5 => UNWINDOWED_174 ,
										MUX_10_1_IN_6 => UNWINDOWED_174 ,
										MUX_10_1_IN_7 => UNWINDOWED_47 ,
										MUX_10_1_IN_8 => UNWINDOWED_302 ,
										MUX_10_1_IN_9 => UNWINDOWED_302 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_151
									);
MUX_REORD_UNIT_152 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_152 ,
										MUX_10_1_IN_1 => UNWINDOWED_152 ,
										MUX_10_1_IN_2 => UNWINDOWED_152 ,
										MUX_10_1_IN_3 => UNWINDOWED_145 ,
										MUX_10_1_IN_4 => UNWINDOWED_145 ,
										MUX_10_1_IN_5 => UNWINDOWED_176 ,
										MUX_10_1_IN_6 => UNWINDOWED_176 ,
										MUX_10_1_IN_7 => UNWINDOWED_49 ,
										MUX_10_1_IN_8 => UNWINDOWED_304 ,
										MUX_10_1_IN_9 => UNWINDOWED_304 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_152
									);
MUX_REORD_UNIT_153 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_153 ,
										MUX_10_1_IN_1 => UNWINDOWED_154 ,
										MUX_10_1_IN_2 => UNWINDOWED_154 ,
										MUX_10_1_IN_3 => UNWINDOWED_147 ,
										MUX_10_1_IN_4 => UNWINDOWED_147 ,
										MUX_10_1_IN_5 => UNWINDOWED_178 ,
										MUX_10_1_IN_6 => UNWINDOWED_178 ,
										MUX_10_1_IN_7 => UNWINDOWED_51 ,
										MUX_10_1_IN_8 => UNWINDOWED_306 ,
										MUX_10_1_IN_9 => UNWINDOWED_306 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_153
									);
MUX_REORD_UNIT_154 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_154 ,
										MUX_10_1_IN_1 => UNWINDOWED_153 ,
										MUX_10_1_IN_2 => UNWINDOWED_156 ,
										MUX_10_1_IN_3 => UNWINDOWED_149 ,
										MUX_10_1_IN_4 => UNWINDOWED_149 ,
										MUX_10_1_IN_5 => UNWINDOWED_180 ,
										MUX_10_1_IN_6 => UNWINDOWED_180 ,
										MUX_10_1_IN_7 => UNWINDOWED_53 ,
										MUX_10_1_IN_8 => UNWINDOWED_308 ,
										MUX_10_1_IN_9 => UNWINDOWED_308 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_154
									);
MUX_REORD_UNIT_155 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_155 ,
										MUX_10_1_IN_1 => UNWINDOWED_155 ,
										MUX_10_1_IN_2 => UNWINDOWED_158 ,
										MUX_10_1_IN_3 => UNWINDOWED_151 ,
										MUX_10_1_IN_4 => UNWINDOWED_151 ,
										MUX_10_1_IN_5 => UNWINDOWED_182 ,
										MUX_10_1_IN_6 => UNWINDOWED_182 ,
										MUX_10_1_IN_7 => UNWINDOWED_55 ,
										MUX_10_1_IN_8 => UNWINDOWED_310 ,
										MUX_10_1_IN_9 => UNWINDOWED_310 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_155
									);
MUX_REORD_UNIT_156 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_156 ,
										MUX_10_1_IN_1 => UNWINDOWED_156 ,
										MUX_10_1_IN_2 => UNWINDOWED_153 ,
										MUX_10_1_IN_3 => UNWINDOWED_153 ,
										MUX_10_1_IN_4 => UNWINDOWED_153 ,
										MUX_10_1_IN_5 => UNWINDOWED_184 ,
										MUX_10_1_IN_6 => UNWINDOWED_184 ,
										MUX_10_1_IN_7 => UNWINDOWED_57 ,
										MUX_10_1_IN_8 => UNWINDOWED_312 ,
										MUX_10_1_IN_9 => UNWINDOWED_312 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_156
									);
MUX_REORD_UNIT_157 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_157 ,
										MUX_10_1_IN_1 => UNWINDOWED_158 ,
										MUX_10_1_IN_2 => UNWINDOWED_155 ,
										MUX_10_1_IN_3 => UNWINDOWED_155 ,
										MUX_10_1_IN_4 => UNWINDOWED_155 ,
										MUX_10_1_IN_5 => UNWINDOWED_186 ,
										MUX_10_1_IN_6 => UNWINDOWED_186 ,
										MUX_10_1_IN_7 => UNWINDOWED_59 ,
										MUX_10_1_IN_8 => UNWINDOWED_314 ,
										MUX_10_1_IN_9 => UNWINDOWED_314 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_157
									);
MUX_REORD_UNIT_158 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_158 ,
										MUX_10_1_IN_1 => UNWINDOWED_157 ,
										MUX_10_1_IN_2 => UNWINDOWED_157 ,
										MUX_10_1_IN_3 => UNWINDOWED_157 ,
										MUX_10_1_IN_4 => UNWINDOWED_157 ,
										MUX_10_1_IN_5 => UNWINDOWED_188 ,
										MUX_10_1_IN_6 => UNWINDOWED_188 ,
										MUX_10_1_IN_7 => UNWINDOWED_61 ,
										MUX_10_1_IN_8 => UNWINDOWED_316 ,
										MUX_10_1_IN_9 => UNWINDOWED_316 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_158
									);
MUX_REORD_UNIT_159 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_159 ,
										MUX_10_1_IN_1 => UNWINDOWED_159 ,
										MUX_10_1_IN_2 => UNWINDOWED_159 ,
										MUX_10_1_IN_3 => UNWINDOWED_159 ,
										MUX_10_1_IN_4 => UNWINDOWED_159 ,
										MUX_10_1_IN_5 => UNWINDOWED_190 ,
										MUX_10_1_IN_6 => UNWINDOWED_190 ,
										MUX_10_1_IN_7 => UNWINDOWED_63 ,
										MUX_10_1_IN_8 => UNWINDOWED_318 ,
										MUX_10_1_IN_9 => UNWINDOWED_318 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_159
									);
MUX_REORD_UNIT_160 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_160 ,
										MUX_10_1_IN_1 => UNWINDOWED_160 ,
										MUX_10_1_IN_2 => UNWINDOWED_160 ,
										MUX_10_1_IN_3 => UNWINDOWED_160 ,
										MUX_10_1_IN_4 => UNWINDOWED_160 ,
										MUX_10_1_IN_5 => UNWINDOWED_129 ,
										MUX_10_1_IN_6 => UNWINDOWED_192 ,
										MUX_10_1_IN_7 => UNWINDOWED_65 ,
										MUX_10_1_IN_8 => UNWINDOWED_320 ,
										MUX_10_1_IN_9 => UNWINDOWED_320 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_160
									);
MUX_REORD_UNIT_161 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_161 ,
										MUX_10_1_IN_1 => UNWINDOWED_162 ,
										MUX_10_1_IN_2 => UNWINDOWED_162 ,
										MUX_10_1_IN_3 => UNWINDOWED_162 ,
										MUX_10_1_IN_4 => UNWINDOWED_162 ,
										MUX_10_1_IN_5 => UNWINDOWED_131 ,
										MUX_10_1_IN_6 => UNWINDOWED_194 ,
										MUX_10_1_IN_7 => UNWINDOWED_67 ,
										MUX_10_1_IN_8 => UNWINDOWED_322 ,
										MUX_10_1_IN_9 => UNWINDOWED_322 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_161
									);
MUX_REORD_UNIT_162 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_162 ,
										MUX_10_1_IN_1 => UNWINDOWED_161 ,
										MUX_10_1_IN_2 => UNWINDOWED_164 ,
										MUX_10_1_IN_3 => UNWINDOWED_164 ,
										MUX_10_1_IN_4 => UNWINDOWED_164 ,
										MUX_10_1_IN_5 => UNWINDOWED_133 ,
										MUX_10_1_IN_6 => UNWINDOWED_196 ,
										MUX_10_1_IN_7 => UNWINDOWED_69 ,
										MUX_10_1_IN_8 => UNWINDOWED_324 ,
										MUX_10_1_IN_9 => UNWINDOWED_324 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_162
									);
MUX_REORD_UNIT_163 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_163 ,
										MUX_10_1_IN_1 => UNWINDOWED_163 ,
										MUX_10_1_IN_2 => UNWINDOWED_166 ,
										MUX_10_1_IN_3 => UNWINDOWED_166 ,
										MUX_10_1_IN_4 => UNWINDOWED_166 ,
										MUX_10_1_IN_5 => UNWINDOWED_135 ,
										MUX_10_1_IN_6 => UNWINDOWED_198 ,
										MUX_10_1_IN_7 => UNWINDOWED_71 ,
										MUX_10_1_IN_8 => UNWINDOWED_326 ,
										MUX_10_1_IN_9 => UNWINDOWED_326 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_163
									);
MUX_REORD_UNIT_164 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_164 ,
										MUX_10_1_IN_1 => UNWINDOWED_164 ,
										MUX_10_1_IN_2 => UNWINDOWED_161 ,
										MUX_10_1_IN_3 => UNWINDOWED_168 ,
										MUX_10_1_IN_4 => UNWINDOWED_168 ,
										MUX_10_1_IN_5 => UNWINDOWED_137 ,
										MUX_10_1_IN_6 => UNWINDOWED_200 ,
										MUX_10_1_IN_7 => UNWINDOWED_73 ,
										MUX_10_1_IN_8 => UNWINDOWED_328 ,
										MUX_10_1_IN_9 => UNWINDOWED_328 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_164
									);
MUX_REORD_UNIT_165 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_165 ,
										MUX_10_1_IN_1 => UNWINDOWED_166 ,
										MUX_10_1_IN_2 => UNWINDOWED_163 ,
										MUX_10_1_IN_3 => UNWINDOWED_170 ,
										MUX_10_1_IN_4 => UNWINDOWED_170 ,
										MUX_10_1_IN_5 => UNWINDOWED_139 ,
										MUX_10_1_IN_6 => UNWINDOWED_202 ,
										MUX_10_1_IN_7 => UNWINDOWED_75 ,
										MUX_10_1_IN_8 => UNWINDOWED_330 ,
										MUX_10_1_IN_9 => UNWINDOWED_330 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_165
									);
MUX_REORD_UNIT_166 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_166 ,
										MUX_10_1_IN_1 => UNWINDOWED_165 ,
										MUX_10_1_IN_2 => UNWINDOWED_165 ,
										MUX_10_1_IN_3 => UNWINDOWED_172 ,
										MUX_10_1_IN_4 => UNWINDOWED_172 ,
										MUX_10_1_IN_5 => UNWINDOWED_141 ,
										MUX_10_1_IN_6 => UNWINDOWED_204 ,
										MUX_10_1_IN_7 => UNWINDOWED_77 ,
										MUX_10_1_IN_8 => UNWINDOWED_332 ,
										MUX_10_1_IN_9 => UNWINDOWED_332 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_166
									);
MUX_REORD_UNIT_167 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_167 ,
										MUX_10_1_IN_1 => UNWINDOWED_167 ,
										MUX_10_1_IN_2 => UNWINDOWED_167 ,
										MUX_10_1_IN_3 => UNWINDOWED_174 ,
										MUX_10_1_IN_4 => UNWINDOWED_174 ,
										MUX_10_1_IN_5 => UNWINDOWED_143 ,
										MUX_10_1_IN_6 => UNWINDOWED_206 ,
										MUX_10_1_IN_7 => UNWINDOWED_79 ,
										MUX_10_1_IN_8 => UNWINDOWED_334 ,
										MUX_10_1_IN_9 => UNWINDOWED_334 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_167
									);
MUX_REORD_UNIT_168 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_168 ,
										MUX_10_1_IN_1 => UNWINDOWED_168 ,
										MUX_10_1_IN_2 => UNWINDOWED_168 ,
										MUX_10_1_IN_3 => UNWINDOWED_161 ,
										MUX_10_1_IN_4 => UNWINDOWED_176 ,
										MUX_10_1_IN_5 => UNWINDOWED_145 ,
										MUX_10_1_IN_6 => UNWINDOWED_208 ,
										MUX_10_1_IN_7 => UNWINDOWED_81 ,
										MUX_10_1_IN_8 => UNWINDOWED_336 ,
										MUX_10_1_IN_9 => UNWINDOWED_336 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_168
									);
MUX_REORD_UNIT_169 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_169 ,
										MUX_10_1_IN_1 => UNWINDOWED_170 ,
										MUX_10_1_IN_2 => UNWINDOWED_170 ,
										MUX_10_1_IN_3 => UNWINDOWED_163 ,
										MUX_10_1_IN_4 => UNWINDOWED_178 ,
										MUX_10_1_IN_5 => UNWINDOWED_147 ,
										MUX_10_1_IN_6 => UNWINDOWED_210 ,
										MUX_10_1_IN_7 => UNWINDOWED_83 ,
										MUX_10_1_IN_8 => UNWINDOWED_338 ,
										MUX_10_1_IN_9 => UNWINDOWED_338 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_169
									);
MUX_REORD_UNIT_170 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_170 ,
										MUX_10_1_IN_1 => UNWINDOWED_169 ,
										MUX_10_1_IN_2 => UNWINDOWED_172 ,
										MUX_10_1_IN_3 => UNWINDOWED_165 ,
										MUX_10_1_IN_4 => UNWINDOWED_180 ,
										MUX_10_1_IN_5 => UNWINDOWED_149 ,
										MUX_10_1_IN_6 => UNWINDOWED_212 ,
										MUX_10_1_IN_7 => UNWINDOWED_85 ,
										MUX_10_1_IN_8 => UNWINDOWED_340 ,
										MUX_10_1_IN_9 => UNWINDOWED_340 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_170
									);
MUX_REORD_UNIT_171 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_171 ,
										MUX_10_1_IN_1 => UNWINDOWED_171 ,
										MUX_10_1_IN_2 => UNWINDOWED_174 ,
										MUX_10_1_IN_3 => UNWINDOWED_167 ,
										MUX_10_1_IN_4 => UNWINDOWED_182 ,
										MUX_10_1_IN_5 => UNWINDOWED_151 ,
										MUX_10_1_IN_6 => UNWINDOWED_214 ,
										MUX_10_1_IN_7 => UNWINDOWED_87 ,
										MUX_10_1_IN_8 => UNWINDOWED_342 ,
										MUX_10_1_IN_9 => UNWINDOWED_342 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_171
									);
MUX_REORD_UNIT_172 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_172 ,
										MUX_10_1_IN_1 => UNWINDOWED_172 ,
										MUX_10_1_IN_2 => UNWINDOWED_169 ,
										MUX_10_1_IN_3 => UNWINDOWED_169 ,
										MUX_10_1_IN_4 => UNWINDOWED_184 ,
										MUX_10_1_IN_5 => UNWINDOWED_153 ,
										MUX_10_1_IN_6 => UNWINDOWED_216 ,
										MUX_10_1_IN_7 => UNWINDOWED_89 ,
										MUX_10_1_IN_8 => UNWINDOWED_344 ,
										MUX_10_1_IN_9 => UNWINDOWED_344 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_172
									);
MUX_REORD_UNIT_173 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_173 ,
										MUX_10_1_IN_1 => UNWINDOWED_174 ,
										MUX_10_1_IN_2 => UNWINDOWED_171 ,
										MUX_10_1_IN_3 => UNWINDOWED_171 ,
										MUX_10_1_IN_4 => UNWINDOWED_186 ,
										MUX_10_1_IN_5 => UNWINDOWED_155 ,
										MUX_10_1_IN_6 => UNWINDOWED_218 ,
										MUX_10_1_IN_7 => UNWINDOWED_91 ,
										MUX_10_1_IN_8 => UNWINDOWED_346 ,
										MUX_10_1_IN_9 => UNWINDOWED_346 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_173
									);
MUX_REORD_UNIT_174 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_174 ,
										MUX_10_1_IN_1 => UNWINDOWED_173 ,
										MUX_10_1_IN_2 => UNWINDOWED_173 ,
										MUX_10_1_IN_3 => UNWINDOWED_173 ,
										MUX_10_1_IN_4 => UNWINDOWED_188 ,
										MUX_10_1_IN_5 => UNWINDOWED_157 ,
										MUX_10_1_IN_6 => UNWINDOWED_220 ,
										MUX_10_1_IN_7 => UNWINDOWED_93 ,
										MUX_10_1_IN_8 => UNWINDOWED_348 ,
										MUX_10_1_IN_9 => UNWINDOWED_348 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_174
									);
MUX_REORD_UNIT_175 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_175 ,
										MUX_10_1_IN_1 => UNWINDOWED_175 ,
										MUX_10_1_IN_2 => UNWINDOWED_175 ,
										MUX_10_1_IN_3 => UNWINDOWED_175 ,
										MUX_10_1_IN_4 => UNWINDOWED_190 ,
										MUX_10_1_IN_5 => UNWINDOWED_159 ,
										MUX_10_1_IN_6 => UNWINDOWED_222 ,
										MUX_10_1_IN_7 => UNWINDOWED_95 ,
										MUX_10_1_IN_8 => UNWINDOWED_350 ,
										MUX_10_1_IN_9 => UNWINDOWED_350 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_175
									);
MUX_REORD_UNIT_176 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_176 ,
										MUX_10_1_IN_1 => UNWINDOWED_176 ,
										MUX_10_1_IN_2 => UNWINDOWED_176 ,
										MUX_10_1_IN_3 => UNWINDOWED_176 ,
										MUX_10_1_IN_4 => UNWINDOWED_161 ,
										MUX_10_1_IN_5 => UNWINDOWED_161 ,
										MUX_10_1_IN_6 => UNWINDOWED_224 ,
										MUX_10_1_IN_7 => UNWINDOWED_97 ,
										MUX_10_1_IN_8 => UNWINDOWED_352 ,
										MUX_10_1_IN_9 => UNWINDOWED_352 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_176
									);
MUX_REORD_UNIT_177 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_177 ,
										MUX_10_1_IN_1 => UNWINDOWED_178 ,
										MUX_10_1_IN_2 => UNWINDOWED_178 ,
										MUX_10_1_IN_3 => UNWINDOWED_178 ,
										MUX_10_1_IN_4 => UNWINDOWED_163 ,
										MUX_10_1_IN_5 => UNWINDOWED_163 ,
										MUX_10_1_IN_6 => UNWINDOWED_226 ,
										MUX_10_1_IN_7 => UNWINDOWED_99 ,
										MUX_10_1_IN_8 => UNWINDOWED_354 ,
										MUX_10_1_IN_9 => UNWINDOWED_354 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_177
									);
MUX_REORD_UNIT_178 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_178 ,
										MUX_10_1_IN_1 => UNWINDOWED_177 ,
										MUX_10_1_IN_2 => UNWINDOWED_180 ,
										MUX_10_1_IN_3 => UNWINDOWED_180 ,
										MUX_10_1_IN_4 => UNWINDOWED_165 ,
										MUX_10_1_IN_5 => UNWINDOWED_165 ,
										MUX_10_1_IN_6 => UNWINDOWED_228 ,
										MUX_10_1_IN_7 => UNWINDOWED_101 ,
										MUX_10_1_IN_8 => UNWINDOWED_356 ,
										MUX_10_1_IN_9 => UNWINDOWED_356 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_178
									);
MUX_REORD_UNIT_179 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_179 ,
										MUX_10_1_IN_1 => UNWINDOWED_179 ,
										MUX_10_1_IN_2 => UNWINDOWED_182 ,
										MUX_10_1_IN_3 => UNWINDOWED_182 ,
										MUX_10_1_IN_4 => UNWINDOWED_167 ,
										MUX_10_1_IN_5 => UNWINDOWED_167 ,
										MUX_10_1_IN_6 => UNWINDOWED_230 ,
										MUX_10_1_IN_7 => UNWINDOWED_103 ,
										MUX_10_1_IN_8 => UNWINDOWED_358 ,
										MUX_10_1_IN_9 => UNWINDOWED_358 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_179
									);
MUX_REORD_UNIT_180 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_180 ,
										MUX_10_1_IN_1 => UNWINDOWED_180 ,
										MUX_10_1_IN_2 => UNWINDOWED_177 ,
										MUX_10_1_IN_3 => UNWINDOWED_184 ,
										MUX_10_1_IN_4 => UNWINDOWED_169 ,
										MUX_10_1_IN_5 => UNWINDOWED_169 ,
										MUX_10_1_IN_6 => UNWINDOWED_232 ,
										MUX_10_1_IN_7 => UNWINDOWED_105 ,
										MUX_10_1_IN_8 => UNWINDOWED_360 ,
										MUX_10_1_IN_9 => UNWINDOWED_360 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_180
									);
MUX_REORD_UNIT_181 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_181 ,
										MUX_10_1_IN_1 => UNWINDOWED_182 ,
										MUX_10_1_IN_2 => UNWINDOWED_179 ,
										MUX_10_1_IN_3 => UNWINDOWED_186 ,
										MUX_10_1_IN_4 => UNWINDOWED_171 ,
										MUX_10_1_IN_5 => UNWINDOWED_171 ,
										MUX_10_1_IN_6 => UNWINDOWED_234 ,
										MUX_10_1_IN_7 => UNWINDOWED_107 ,
										MUX_10_1_IN_8 => UNWINDOWED_362 ,
										MUX_10_1_IN_9 => UNWINDOWED_362 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_181
									);
MUX_REORD_UNIT_182 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_182 ,
										MUX_10_1_IN_1 => UNWINDOWED_181 ,
										MUX_10_1_IN_2 => UNWINDOWED_181 ,
										MUX_10_1_IN_3 => UNWINDOWED_188 ,
										MUX_10_1_IN_4 => UNWINDOWED_173 ,
										MUX_10_1_IN_5 => UNWINDOWED_173 ,
										MUX_10_1_IN_6 => UNWINDOWED_236 ,
										MUX_10_1_IN_7 => UNWINDOWED_109 ,
										MUX_10_1_IN_8 => UNWINDOWED_364 ,
										MUX_10_1_IN_9 => UNWINDOWED_364 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_182
									);
MUX_REORD_UNIT_183 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_183 ,
										MUX_10_1_IN_1 => UNWINDOWED_183 ,
										MUX_10_1_IN_2 => UNWINDOWED_183 ,
										MUX_10_1_IN_3 => UNWINDOWED_190 ,
										MUX_10_1_IN_4 => UNWINDOWED_175 ,
										MUX_10_1_IN_5 => UNWINDOWED_175 ,
										MUX_10_1_IN_6 => UNWINDOWED_238 ,
										MUX_10_1_IN_7 => UNWINDOWED_111 ,
										MUX_10_1_IN_8 => UNWINDOWED_366 ,
										MUX_10_1_IN_9 => UNWINDOWED_366 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_183
									);
MUX_REORD_UNIT_184 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_184 ,
										MUX_10_1_IN_1 => UNWINDOWED_184 ,
										MUX_10_1_IN_2 => UNWINDOWED_184 ,
										MUX_10_1_IN_3 => UNWINDOWED_177 ,
										MUX_10_1_IN_4 => UNWINDOWED_177 ,
										MUX_10_1_IN_5 => UNWINDOWED_177 ,
										MUX_10_1_IN_6 => UNWINDOWED_240 ,
										MUX_10_1_IN_7 => UNWINDOWED_113 ,
										MUX_10_1_IN_8 => UNWINDOWED_368 ,
										MUX_10_1_IN_9 => UNWINDOWED_368 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_184
									);
MUX_REORD_UNIT_185 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_185 ,
										MUX_10_1_IN_1 => UNWINDOWED_186 ,
										MUX_10_1_IN_2 => UNWINDOWED_186 ,
										MUX_10_1_IN_3 => UNWINDOWED_179 ,
										MUX_10_1_IN_4 => UNWINDOWED_179 ,
										MUX_10_1_IN_5 => UNWINDOWED_179 ,
										MUX_10_1_IN_6 => UNWINDOWED_242 ,
										MUX_10_1_IN_7 => UNWINDOWED_115 ,
										MUX_10_1_IN_8 => UNWINDOWED_370 ,
										MUX_10_1_IN_9 => UNWINDOWED_370 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_185
									);
MUX_REORD_UNIT_186 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_186 ,
										MUX_10_1_IN_1 => UNWINDOWED_185 ,
										MUX_10_1_IN_2 => UNWINDOWED_188 ,
										MUX_10_1_IN_3 => UNWINDOWED_181 ,
										MUX_10_1_IN_4 => UNWINDOWED_181 ,
										MUX_10_1_IN_5 => UNWINDOWED_181 ,
										MUX_10_1_IN_6 => UNWINDOWED_244 ,
										MUX_10_1_IN_7 => UNWINDOWED_117 ,
										MUX_10_1_IN_8 => UNWINDOWED_372 ,
										MUX_10_1_IN_9 => UNWINDOWED_372 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_186
									);
MUX_REORD_UNIT_187 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_187 ,
										MUX_10_1_IN_1 => UNWINDOWED_187 ,
										MUX_10_1_IN_2 => UNWINDOWED_190 ,
										MUX_10_1_IN_3 => UNWINDOWED_183 ,
										MUX_10_1_IN_4 => UNWINDOWED_183 ,
										MUX_10_1_IN_5 => UNWINDOWED_183 ,
										MUX_10_1_IN_6 => UNWINDOWED_246 ,
										MUX_10_1_IN_7 => UNWINDOWED_119 ,
										MUX_10_1_IN_8 => UNWINDOWED_374 ,
										MUX_10_1_IN_9 => UNWINDOWED_374 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_187
									);
MUX_REORD_UNIT_188 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_188 ,
										MUX_10_1_IN_1 => UNWINDOWED_188 ,
										MUX_10_1_IN_2 => UNWINDOWED_185 ,
										MUX_10_1_IN_3 => UNWINDOWED_185 ,
										MUX_10_1_IN_4 => UNWINDOWED_185 ,
										MUX_10_1_IN_5 => UNWINDOWED_185 ,
										MUX_10_1_IN_6 => UNWINDOWED_248 ,
										MUX_10_1_IN_7 => UNWINDOWED_121 ,
										MUX_10_1_IN_8 => UNWINDOWED_376 ,
										MUX_10_1_IN_9 => UNWINDOWED_376 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_188
									);
MUX_REORD_UNIT_189 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_189 ,
										MUX_10_1_IN_1 => UNWINDOWED_190 ,
										MUX_10_1_IN_2 => UNWINDOWED_187 ,
										MUX_10_1_IN_3 => UNWINDOWED_187 ,
										MUX_10_1_IN_4 => UNWINDOWED_187 ,
										MUX_10_1_IN_5 => UNWINDOWED_187 ,
										MUX_10_1_IN_6 => UNWINDOWED_250 ,
										MUX_10_1_IN_7 => UNWINDOWED_123 ,
										MUX_10_1_IN_8 => UNWINDOWED_378 ,
										MUX_10_1_IN_9 => UNWINDOWED_378 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_189
									);
MUX_REORD_UNIT_190 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_190 ,
										MUX_10_1_IN_1 => UNWINDOWED_189 ,
										MUX_10_1_IN_2 => UNWINDOWED_189 ,
										MUX_10_1_IN_3 => UNWINDOWED_189 ,
										MUX_10_1_IN_4 => UNWINDOWED_189 ,
										MUX_10_1_IN_5 => UNWINDOWED_189 ,
										MUX_10_1_IN_6 => UNWINDOWED_252 ,
										MUX_10_1_IN_7 => UNWINDOWED_125 ,
										MUX_10_1_IN_8 => UNWINDOWED_380 ,
										MUX_10_1_IN_9 => UNWINDOWED_380 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_190
									);
MUX_REORD_UNIT_191 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_191 ,
										MUX_10_1_IN_1 => UNWINDOWED_191 ,
										MUX_10_1_IN_2 => UNWINDOWED_191 ,
										MUX_10_1_IN_3 => UNWINDOWED_191 ,
										MUX_10_1_IN_4 => UNWINDOWED_191 ,
										MUX_10_1_IN_5 => UNWINDOWED_191 ,
										MUX_10_1_IN_6 => UNWINDOWED_254 ,
										MUX_10_1_IN_7 => UNWINDOWED_127 ,
										MUX_10_1_IN_8 => UNWINDOWED_382 ,
										MUX_10_1_IN_9 => UNWINDOWED_382 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_191
									);
MUX_REORD_UNIT_192 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_192 ,
										MUX_10_1_IN_1 => UNWINDOWED_192 ,
										MUX_10_1_IN_2 => UNWINDOWED_192 ,
										MUX_10_1_IN_3 => UNWINDOWED_192 ,
										MUX_10_1_IN_4 => UNWINDOWED_192 ,
										MUX_10_1_IN_5 => UNWINDOWED_192 ,
										MUX_10_1_IN_6 => UNWINDOWED_129 ,
										MUX_10_1_IN_7 => UNWINDOWED_129 ,
										MUX_10_1_IN_8 => UNWINDOWED_384 ,
										MUX_10_1_IN_9 => UNWINDOWED_384 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_192
									);
MUX_REORD_UNIT_193 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_193 ,
										MUX_10_1_IN_1 => UNWINDOWED_194 ,
										MUX_10_1_IN_2 => UNWINDOWED_194 ,
										MUX_10_1_IN_3 => UNWINDOWED_194 ,
										MUX_10_1_IN_4 => UNWINDOWED_194 ,
										MUX_10_1_IN_5 => UNWINDOWED_194 ,
										MUX_10_1_IN_6 => UNWINDOWED_131 ,
										MUX_10_1_IN_7 => UNWINDOWED_131 ,
										MUX_10_1_IN_8 => UNWINDOWED_386 ,
										MUX_10_1_IN_9 => UNWINDOWED_386 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_193
									);
MUX_REORD_UNIT_194 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_194 ,
										MUX_10_1_IN_1 => UNWINDOWED_193 ,
										MUX_10_1_IN_2 => UNWINDOWED_196 ,
										MUX_10_1_IN_3 => UNWINDOWED_196 ,
										MUX_10_1_IN_4 => UNWINDOWED_196 ,
										MUX_10_1_IN_5 => UNWINDOWED_196 ,
										MUX_10_1_IN_6 => UNWINDOWED_133 ,
										MUX_10_1_IN_7 => UNWINDOWED_133 ,
										MUX_10_1_IN_8 => UNWINDOWED_388 ,
										MUX_10_1_IN_9 => UNWINDOWED_388 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_194
									);
MUX_REORD_UNIT_195 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_195 ,
										MUX_10_1_IN_1 => UNWINDOWED_195 ,
										MUX_10_1_IN_2 => UNWINDOWED_198 ,
										MUX_10_1_IN_3 => UNWINDOWED_198 ,
										MUX_10_1_IN_4 => UNWINDOWED_198 ,
										MUX_10_1_IN_5 => UNWINDOWED_198 ,
										MUX_10_1_IN_6 => UNWINDOWED_135 ,
										MUX_10_1_IN_7 => UNWINDOWED_135 ,
										MUX_10_1_IN_8 => UNWINDOWED_390 ,
										MUX_10_1_IN_9 => UNWINDOWED_390 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_195
									);
MUX_REORD_UNIT_196 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_196 ,
										MUX_10_1_IN_1 => UNWINDOWED_196 ,
										MUX_10_1_IN_2 => UNWINDOWED_193 ,
										MUX_10_1_IN_3 => UNWINDOWED_200 ,
										MUX_10_1_IN_4 => UNWINDOWED_200 ,
										MUX_10_1_IN_5 => UNWINDOWED_200 ,
										MUX_10_1_IN_6 => UNWINDOWED_137 ,
										MUX_10_1_IN_7 => UNWINDOWED_137 ,
										MUX_10_1_IN_8 => UNWINDOWED_392 ,
										MUX_10_1_IN_9 => UNWINDOWED_392 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_196
									);
MUX_REORD_UNIT_197 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_197 ,
										MUX_10_1_IN_1 => UNWINDOWED_198 ,
										MUX_10_1_IN_2 => UNWINDOWED_195 ,
										MUX_10_1_IN_3 => UNWINDOWED_202 ,
										MUX_10_1_IN_4 => UNWINDOWED_202 ,
										MUX_10_1_IN_5 => UNWINDOWED_202 ,
										MUX_10_1_IN_6 => UNWINDOWED_139 ,
										MUX_10_1_IN_7 => UNWINDOWED_139 ,
										MUX_10_1_IN_8 => UNWINDOWED_394 ,
										MUX_10_1_IN_9 => UNWINDOWED_394 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_197
									);
MUX_REORD_UNIT_198 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_198 ,
										MUX_10_1_IN_1 => UNWINDOWED_197 ,
										MUX_10_1_IN_2 => UNWINDOWED_197 ,
										MUX_10_1_IN_3 => UNWINDOWED_204 ,
										MUX_10_1_IN_4 => UNWINDOWED_204 ,
										MUX_10_1_IN_5 => UNWINDOWED_204 ,
										MUX_10_1_IN_6 => UNWINDOWED_141 ,
										MUX_10_1_IN_7 => UNWINDOWED_141 ,
										MUX_10_1_IN_8 => UNWINDOWED_396 ,
										MUX_10_1_IN_9 => UNWINDOWED_396 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_198
									);
MUX_REORD_UNIT_199 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_199 ,
										MUX_10_1_IN_1 => UNWINDOWED_199 ,
										MUX_10_1_IN_2 => UNWINDOWED_199 ,
										MUX_10_1_IN_3 => UNWINDOWED_206 ,
										MUX_10_1_IN_4 => UNWINDOWED_206 ,
										MUX_10_1_IN_5 => UNWINDOWED_206 ,
										MUX_10_1_IN_6 => UNWINDOWED_143 ,
										MUX_10_1_IN_7 => UNWINDOWED_143 ,
										MUX_10_1_IN_8 => UNWINDOWED_398 ,
										MUX_10_1_IN_9 => UNWINDOWED_398 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_199
									);
MUX_REORD_UNIT_200 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_200 ,
										MUX_10_1_IN_1 => UNWINDOWED_200 ,
										MUX_10_1_IN_2 => UNWINDOWED_200 ,
										MUX_10_1_IN_3 => UNWINDOWED_193 ,
										MUX_10_1_IN_4 => UNWINDOWED_208 ,
										MUX_10_1_IN_5 => UNWINDOWED_208 ,
										MUX_10_1_IN_6 => UNWINDOWED_145 ,
										MUX_10_1_IN_7 => UNWINDOWED_145 ,
										MUX_10_1_IN_8 => UNWINDOWED_400 ,
										MUX_10_1_IN_9 => UNWINDOWED_400 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_200
									);
MUX_REORD_UNIT_201 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_201 ,
										MUX_10_1_IN_1 => UNWINDOWED_202 ,
										MUX_10_1_IN_2 => UNWINDOWED_202 ,
										MUX_10_1_IN_3 => UNWINDOWED_195 ,
										MUX_10_1_IN_4 => UNWINDOWED_210 ,
										MUX_10_1_IN_5 => UNWINDOWED_210 ,
										MUX_10_1_IN_6 => UNWINDOWED_147 ,
										MUX_10_1_IN_7 => UNWINDOWED_147 ,
										MUX_10_1_IN_8 => UNWINDOWED_402 ,
										MUX_10_1_IN_9 => UNWINDOWED_402 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_201
									);
MUX_REORD_UNIT_202 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_202 ,
										MUX_10_1_IN_1 => UNWINDOWED_201 ,
										MUX_10_1_IN_2 => UNWINDOWED_204 ,
										MUX_10_1_IN_3 => UNWINDOWED_197 ,
										MUX_10_1_IN_4 => UNWINDOWED_212 ,
										MUX_10_1_IN_5 => UNWINDOWED_212 ,
										MUX_10_1_IN_6 => UNWINDOWED_149 ,
										MUX_10_1_IN_7 => UNWINDOWED_149 ,
										MUX_10_1_IN_8 => UNWINDOWED_404 ,
										MUX_10_1_IN_9 => UNWINDOWED_404 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_202
									);
MUX_REORD_UNIT_203 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_203 ,
										MUX_10_1_IN_1 => UNWINDOWED_203 ,
										MUX_10_1_IN_2 => UNWINDOWED_206 ,
										MUX_10_1_IN_3 => UNWINDOWED_199 ,
										MUX_10_1_IN_4 => UNWINDOWED_214 ,
										MUX_10_1_IN_5 => UNWINDOWED_214 ,
										MUX_10_1_IN_6 => UNWINDOWED_151 ,
										MUX_10_1_IN_7 => UNWINDOWED_151 ,
										MUX_10_1_IN_8 => UNWINDOWED_406 ,
										MUX_10_1_IN_9 => UNWINDOWED_406 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_203
									);
MUX_REORD_UNIT_204 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_204 ,
										MUX_10_1_IN_1 => UNWINDOWED_204 ,
										MUX_10_1_IN_2 => UNWINDOWED_201 ,
										MUX_10_1_IN_3 => UNWINDOWED_201 ,
										MUX_10_1_IN_4 => UNWINDOWED_216 ,
										MUX_10_1_IN_5 => UNWINDOWED_216 ,
										MUX_10_1_IN_6 => UNWINDOWED_153 ,
										MUX_10_1_IN_7 => UNWINDOWED_153 ,
										MUX_10_1_IN_8 => UNWINDOWED_408 ,
										MUX_10_1_IN_9 => UNWINDOWED_408 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_204
									);
MUX_REORD_UNIT_205 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_205 ,
										MUX_10_1_IN_1 => UNWINDOWED_206 ,
										MUX_10_1_IN_2 => UNWINDOWED_203 ,
										MUX_10_1_IN_3 => UNWINDOWED_203 ,
										MUX_10_1_IN_4 => UNWINDOWED_218 ,
										MUX_10_1_IN_5 => UNWINDOWED_218 ,
										MUX_10_1_IN_6 => UNWINDOWED_155 ,
										MUX_10_1_IN_7 => UNWINDOWED_155 ,
										MUX_10_1_IN_8 => UNWINDOWED_410 ,
										MUX_10_1_IN_9 => UNWINDOWED_410 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_205
									);
MUX_REORD_UNIT_206 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_206 ,
										MUX_10_1_IN_1 => UNWINDOWED_205 ,
										MUX_10_1_IN_2 => UNWINDOWED_205 ,
										MUX_10_1_IN_3 => UNWINDOWED_205 ,
										MUX_10_1_IN_4 => UNWINDOWED_220 ,
										MUX_10_1_IN_5 => UNWINDOWED_220 ,
										MUX_10_1_IN_6 => UNWINDOWED_157 ,
										MUX_10_1_IN_7 => UNWINDOWED_157 ,
										MUX_10_1_IN_8 => UNWINDOWED_412 ,
										MUX_10_1_IN_9 => UNWINDOWED_412 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_206
									);
MUX_REORD_UNIT_207 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_207 ,
										MUX_10_1_IN_1 => UNWINDOWED_207 ,
										MUX_10_1_IN_2 => UNWINDOWED_207 ,
										MUX_10_1_IN_3 => UNWINDOWED_207 ,
										MUX_10_1_IN_4 => UNWINDOWED_222 ,
										MUX_10_1_IN_5 => UNWINDOWED_222 ,
										MUX_10_1_IN_6 => UNWINDOWED_159 ,
										MUX_10_1_IN_7 => UNWINDOWED_159 ,
										MUX_10_1_IN_8 => UNWINDOWED_414 ,
										MUX_10_1_IN_9 => UNWINDOWED_414 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_207
									);
MUX_REORD_UNIT_208 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_208 ,
										MUX_10_1_IN_1 => UNWINDOWED_208 ,
										MUX_10_1_IN_2 => UNWINDOWED_208 ,
										MUX_10_1_IN_3 => UNWINDOWED_208 ,
										MUX_10_1_IN_4 => UNWINDOWED_193 ,
										MUX_10_1_IN_5 => UNWINDOWED_224 ,
										MUX_10_1_IN_6 => UNWINDOWED_161 ,
										MUX_10_1_IN_7 => UNWINDOWED_161 ,
										MUX_10_1_IN_8 => UNWINDOWED_416 ,
										MUX_10_1_IN_9 => UNWINDOWED_416 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_208
									);
MUX_REORD_UNIT_209 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_209 ,
										MUX_10_1_IN_1 => UNWINDOWED_210 ,
										MUX_10_1_IN_2 => UNWINDOWED_210 ,
										MUX_10_1_IN_3 => UNWINDOWED_210 ,
										MUX_10_1_IN_4 => UNWINDOWED_195 ,
										MUX_10_1_IN_5 => UNWINDOWED_226 ,
										MUX_10_1_IN_6 => UNWINDOWED_163 ,
										MUX_10_1_IN_7 => UNWINDOWED_163 ,
										MUX_10_1_IN_8 => UNWINDOWED_418 ,
										MUX_10_1_IN_9 => UNWINDOWED_418 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_209
									);
MUX_REORD_UNIT_210 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_210 ,
										MUX_10_1_IN_1 => UNWINDOWED_209 ,
										MUX_10_1_IN_2 => UNWINDOWED_212 ,
										MUX_10_1_IN_3 => UNWINDOWED_212 ,
										MUX_10_1_IN_4 => UNWINDOWED_197 ,
										MUX_10_1_IN_5 => UNWINDOWED_228 ,
										MUX_10_1_IN_6 => UNWINDOWED_165 ,
										MUX_10_1_IN_7 => UNWINDOWED_165 ,
										MUX_10_1_IN_8 => UNWINDOWED_420 ,
										MUX_10_1_IN_9 => UNWINDOWED_420 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_210
									);
MUX_REORD_UNIT_211 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_211 ,
										MUX_10_1_IN_1 => UNWINDOWED_211 ,
										MUX_10_1_IN_2 => UNWINDOWED_214 ,
										MUX_10_1_IN_3 => UNWINDOWED_214 ,
										MUX_10_1_IN_4 => UNWINDOWED_199 ,
										MUX_10_1_IN_5 => UNWINDOWED_230 ,
										MUX_10_1_IN_6 => UNWINDOWED_167 ,
										MUX_10_1_IN_7 => UNWINDOWED_167 ,
										MUX_10_1_IN_8 => UNWINDOWED_422 ,
										MUX_10_1_IN_9 => UNWINDOWED_422 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_211
									);
MUX_REORD_UNIT_212 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_212 ,
										MUX_10_1_IN_1 => UNWINDOWED_212 ,
										MUX_10_1_IN_2 => UNWINDOWED_209 ,
										MUX_10_1_IN_3 => UNWINDOWED_216 ,
										MUX_10_1_IN_4 => UNWINDOWED_201 ,
										MUX_10_1_IN_5 => UNWINDOWED_232 ,
										MUX_10_1_IN_6 => UNWINDOWED_169 ,
										MUX_10_1_IN_7 => UNWINDOWED_169 ,
										MUX_10_1_IN_8 => UNWINDOWED_424 ,
										MUX_10_1_IN_9 => UNWINDOWED_424 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_212
									);
MUX_REORD_UNIT_213 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_213 ,
										MUX_10_1_IN_1 => UNWINDOWED_214 ,
										MUX_10_1_IN_2 => UNWINDOWED_211 ,
										MUX_10_1_IN_3 => UNWINDOWED_218 ,
										MUX_10_1_IN_4 => UNWINDOWED_203 ,
										MUX_10_1_IN_5 => UNWINDOWED_234 ,
										MUX_10_1_IN_6 => UNWINDOWED_171 ,
										MUX_10_1_IN_7 => UNWINDOWED_171 ,
										MUX_10_1_IN_8 => UNWINDOWED_426 ,
										MUX_10_1_IN_9 => UNWINDOWED_426 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_213
									);
MUX_REORD_UNIT_214 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_214 ,
										MUX_10_1_IN_1 => UNWINDOWED_213 ,
										MUX_10_1_IN_2 => UNWINDOWED_213 ,
										MUX_10_1_IN_3 => UNWINDOWED_220 ,
										MUX_10_1_IN_4 => UNWINDOWED_205 ,
										MUX_10_1_IN_5 => UNWINDOWED_236 ,
										MUX_10_1_IN_6 => UNWINDOWED_173 ,
										MUX_10_1_IN_7 => UNWINDOWED_173 ,
										MUX_10_1_IN_8 => UNWINDOWED_428 ,
										MUX_10_1_IN_9 => UNWINDOWED_428 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_214
									);
MUX_REORD_UNIT_215 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_215 ,
										MUX_10_1_IN_1 => UNWINDOWED_215 ,
										MUX_10_1_IN_2 => UNWINDOWED_215 ,
										MUX_10_1_IN_3 => UNWINDOWED_222 ,
										MUX_10_1_IN_4 => UNWINDOWED_207 ,
										MUX_10_1_IN_5 => UNWINDOWED_238 ,
										MUX_10_1_IN_6 => UNWINDOWED_175 ,
										MUX_10_1_IN_7 => UNWINDOWED_175 ,
										MUX_10_1_IN_8 => UNWINDOWED_430 ,
										MUX_10_1_IN_9 => UNWINDOWED_430 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_215
									);
MUX_REORD_UNIT_216 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_216 ,
										MUX_10_1_IN_1 => UNWINDOWED_216 ,
										MUX_10_1_IN_2 => UNWINDOWED_216 ,
										MUX_10_1_IN_3 => UNWINDOWED_209 ,
										MUX_10_1_IN_4 => UNWINDOWED_209 ,
										MUX_10_1_IN_5 => UNWINDOWED_240 ,
										MUX_10_1_IN_6 => UNWINDOWED_177 ,
										MUX_10_1_IN_7 => UNWINDOWED_177 ,
										MUX_10_1_IN_8 => UNWINDOWED_432 ,
										MUX_10_1_IN_9 => UNWINDOWED_432 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_216
									);
MUX_REORD_UNIT_217 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_217 ,
										MUX_10_1_IN_1 => UNWINDOWED_218 ,
										MUX_10_1_IN_2 => UNWINDOWED_218 ,
										MUX_10_1_IN_3 => UNWINDOWED_211 ,
										MUX_10_1_IN_4 => UNWINDOWED_211 ,
										MUX_10_1_IN_5 => UNWINDOWED_242 ,
										MUX_10_1_IN_6 => UNWINDOWED_179 ,
										MUX_10_1_IN_7 => UNWINDOWED_179 ,
										MUX_10_1_IN_8 => UNWINDOWED_434 ,
										MUX_10_1_IN_9 => UNWINDOWED_434 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_217
									);
MUX_REORD_UNIT_218 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_218 ,
										MUX_10_1_IN_1 => UNWINDOWED_217 ,
										MUX_10_1_IN_2 => UNWINDOWED_220 ,
										MUX_10_1_IN_3 => UNWINDOWED_213 ,
										MUX_10_1_IN_4 => UNWINDOWED_213 ,
										MUX_10_1_IN_5 => UNWINDOWED_244 ,
										MUX_10_1_IN_6 => UNWINDOWED_181 ,
										MUX_10_1_IN_7 => UNWINDOWED_181 ,
										MUX_10_1_IN_8 => UNWINDOWED_436 ,
										MUX_10_1_IN_9 => UNWINDOWED_436 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_218
									);
MUX_REORD_UNIT_219 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_219 ,
										MUX_10_1_IN_1 => UNWINDOWED_219 ,
										MUX_10_1_IN_2 => UNWINDOWED_222 ,
										MUX_10_1_IN_3 => UNWINDOWED_215 ,
										MUX_10_1_IN_4 => UNWINDOWED_215 ,
										MUX_10_1_IN_5 => UNWINDOWED_246 ,
										MUX_10_1_IN_6 => UNWINDOWED_183 ,
										MUX_10_1_IN_7 => UNWINDOWED_183 ,
										MUX_10_1_IN_8 => UNWINDOWED_438 ,
										MUX_10_1_IN_9 => UNWINDOWED_438 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_219
									);
MUX_REORD_UNIT_220 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_220 ,
										MUX_10_1_IN_1 => UNWINDOWED_220 ,
										MUX_10_1_IN_2 => UNWINDOWED_217 ,
										MUX_10_1_IN_3 => UNWINDOWED_217 ,
										MUX_10_1_IN_4 => UNWINDOWED_217 ,
										MUX_10_1_IN_5 => UNWINDOWED_248 ,
										MUX_10_1_IN_6 => UNWINDOWED_185 ,
										MUX_10_1_IN_7 => UNWINDOWED_185 ,
										MUX_10_1_IN_8 => UNWINDOWED_440 ,
										MUX_10_1_IN_9 => UNWINDOWED_440 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_220
									);
MUX_REORD_UNIT_221 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_221 ,
										MUX_10_1_IN_1 => UNWINDOWED_222 ,
										MUX_10_1_IN_2 => UNWINDOWED_219 ,
										MUX_10_1_IN_3 => UNWINDOWED_219 ,
										MUX_10_1_IN_4 => UNWINDOWED_219 ,
										MUX_10_1_IN_5 => UNWINDOWED_250 ,
										MUX_10_1_IN_6 => UNWINDOWED_187 ,
										MUX_10_1_IN_7 => UNWINDOWED_187 ,
										MUX_10_1_IN_8 => UNWINDOWED_442 ,
										MUX_10_1_IN_9 => UNWINDOWED_442 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_221
									);
MUX_REORD_UNIT_222 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_222 ,
										MUX_10_1_IN_1 => UNWINDOWED_221 ,
										MUX_10_1_IN_2 => UNWINDOWED_221 ,
										MUX_10_1_IN_3 => UNWINDOWED_221 ,
										MUX_10_1_IN_4 => UNWINDOWED_221 ,
										MUX_10_1_IN_5 => UNWINDOWED_252 ,
										MUX_10_1_IN_6 => UNWINDOWED_189 ,
										MUX_10_1_IN_7 => UNWINDOWED_189 ,
										MUX_10_1_IN_8 => UNWINDOWED_444 ,
										MUX_10_1_IN_9 => UNWINDOWED_444 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_222
									);
MUX_REORD_UNIT_223 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_223 ,
										MUX_10_1_IN_1 => UNWINDOWED_223 ,
										MUX_10_1_IN_2 => UNWINDOWED_223 ,
										MUX_10_1_IN_3 => UNWINDOWED_223 ,
										MUX_10_1_IN_4 => UNWINDOWED_223 ,
										MUX_10_1_IN_5 => UNWINDOWED_254 ,
										MUX_10_1_IN_6 => UNWINDOWED_191 ,
										MUX_10_1_IN_7 => UNWINDOWED_191 ,
										MUX_10_1_IN_8 => UNWINDOWED_446 ,
										MUX_10_1_IN_9 => UNWINDOWED_446 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_223
									);
MUX_REORD_UNIT_224 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_224 ,
										MUX_10_1_IN_1 => UNWINDOWED_224 ,
										MUX_10_1_IN_2 => UNWINDOWED_224 ,
										MUX_10_1_IN_3 => UNWINDOWED_224 ,
										MUX_10_1_IN_4 => UNWINDOWED_224 ,
										MUX_10_1_IN_5 => UNWINDOWED_193 ,
										MUX_10_1_IN_6 => UNWINDOWED_193 ,
										MUX_10_1_IN_7 => UNWINDOWED_193 ,
										MUX_10_1_IN_8 => UNWINDOWED_448 ,
										MUX_10_1_IN_9 => UNWINDOWED_448 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_224
									);
MUX_REORD_UNIT_225 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_225 ,
										MUX_10_1_IN_1 => UNWINDOWED_226 ,
										MUX_10_1_IN_2 => UNWINDOWED_226 ,
										MUX_10_1_IN_3 => UNWINDOWED_226 ,
										MUX_10_1_IN_4 => UNWINDOWED_226 ,
										MUX_10_1_IN_5 => UNWINDOWED_195 ,
										MUX_10_1_IN_6 => UNWINDOWED_195 ,
										MUX_10_1_IN_7 => UNWINDOWED_195 ,
										MUX_10_1_IN_8 => UNWINDOWED_450 ,
										MUX_10_1_IN_9 => UNWINDOWED_450 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_225
									);
MUX_REORD_UNIT_226 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_226 ,
										MUX_10_1_IN_1 => UNWINDOWED_225 ,
										MUX_10_1_IN_2 => UNWINDOWED_228 ,
										MUX_10_1_IN_3 => UNWINDOWED_228 ,
										MUX_10_1_IN_4 => UNWINDOWED_228 ,
										MUX_10_1_IN_5 => UNWINDOWED_197 ,
										MUX_10_1_IN_6 => UNWINDOWED_197 ,
										MUX_10_1_IN_7 => UNWINDOWED_197 ,
										MUX_10_1_IN_8 => UNWINDOWED_452 ,
										MUX_10_1_IN_9 => UNWINDOWED_452 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_226
									);
MUX_REORD_UNIT_227 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_227 ,
										MUX_10_1_IN_1 => UNWINDOWED_227 ,
										MUX_10_1_IN_2 => UNWINDOWED_230 ,
										MUX_10_1_IN_3 => UNWINDOWED_230 ,
										MUX_10_1_IN_4 => UNWINDOWED_230 ,
										MUX_10_1_IN_5 => UNWINDOWED_199 ,
										MUX_10_1_IN_6 => UNWINDOWED_199 ,
										MUX_10_1_IN_7 => UNWINDOWED_199 ,
										MUX_10_1_IN_8 => UNWINDOWED_454 ,
										MUX_10_1_IN_9 => UNWINDOWED_454 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_227
									);
MUX_REORD_UNIT_228 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_228 ,
										MUX_10_1_IN_1 => UNWINDOWED_228 ,
										MUX_10_1_IN_2 => UNWINDOWED_225 ,
										MUX_10_1_IN_3 => UNWINDOWED_232 ,
										MUX_10_1_IN_4 => UNWINDOWED_232 ,
										MUX_10_1_IN_5 => UNWINDOWED_201 ,
										MUX_10_1_IN_6 => UNWINDOWED_201 ,
										MUX_10_1_IN_7 => UNWINDOWED_201 ,
										MUX_10_1_IN_8 => UNWINDOWED_456 ,
										MUX_10_1_IN_9 => UNWINDOWED_456 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_228
									);
MUX_REORD_UNIT_229 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_229 ,
										MUX_10_1_IN_1 => UNWINDOWED_230 ,
										MUX_10_1_IN_2 => UNWINDOWED_227 ,
										MUX_10_1_IN_3 => UNWINDOWED_234 ,
										MUX_10_1_IN_4 => UNWINDOWED_234 ,
										MUX_10_1_IN_5 => UNWINDOWED_203 ,
										MUX_10_1_IN_6 => UNWINDOWED_203 ,
										MUX_10_1_IN_7 => UNWINDOWED_203 ,
										MUX_10_1_IN_8 => UNWINDOWED_458 ,
										MUX_10_1_IN_9 => UNWINDOWED_458 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_229
									);
MUX_REORD_UNIT_230 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_230 ,
										MUX_10_1_IN_1 => UNWINDOWED_229 ,
										MUX_10_1_IN_2 => UNWINDOWED_229 ,
										MUX_10_1_IN_3 => UNWINDOWED_236 ,
										MUX_10_1_IN_4 => UNWINDOWED_236 ,
										MUX_10_1_IN_5 => UNWINDOWED_205 ,
										MUX_10_1_IN_6 => UNWINDOWED_205 ,
										MUX_10_1_IN_7 => UNWINDOWED_205 ,
										MUX_10_1_IN_8 => UNWINDOWED_460 ,
										MUX_10_1_IN_9 => UNWINDOWED_460 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_230
									);
MUX_REORD_UNIT_231 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_231 ,
										MUX_10_1_IN_1 => UNWINDOWED_231 ,
										MUX_10_1_IN_2 => UNWINDOWED_231 ,
										MUX_10_1_IN_3 => UNWINDOWED_238 ,
										MUX_10_1_IN_4 => UNWINDOWED_238 ,
										MUX_10_1_IN_5 => UNWINDOWED_207 ,
										MUX_10_1_IN_6 => UNWINDOWED_207 ,
										MUX_10_1_IN_7 => UNWINDOWED_207 ,
										MUX_10_1_IN_8 => UNWINDOWED_462 ,
										MUX_10_1_IN_9 => UNWINDOWED_462 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_231
									);
MUX_REORD_UNIT_232 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_232 ,
										MUX_10_1_IN_1 => UNWINDOWED_232 ,
										MUX_10_1_IN_2 => UNWINDOWED_232 ,
										MUX_10_1_IN_3 => UNWINDOWED_225 ,
										MUX_10_1_IN_4 => UNWINDOWED_240 ,
										MUX_10_1_IN_5 => UNWINDOWED_209 ,
										MUX_10_1_IN_6 => UNWINDOWED_209 ,
										MUX_10_1_IN_7 => UNWINDOWED_209 ,
										MUX_10_1_IN_8 => UNWINDOWED_464 ,
										MUX_10_1_IN_9 => UNWINDOWED_464 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_232
									);
MUX_REORD_UNIT_233 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_233 ,
										MUX_10_1_IN_1 => UNWINDOWED_234 ,
										MUX_10_1_IN_2 => UNWINDOWED_234 ,
										MUX_10_1_IN_3 => UNWINDOWED_227 ,
										MUX_10_1_IN_4 => UNWINDOWED_242 ,
										MUX_10_1_IN_5 => UNWINDOWED_211 ,
										MUX_10_1_IN_6 => UNWINDOWED_211 ,
										MUX_10_1_IN_7 => UNWINDOWED_211 ,
										MUX_10_1_IN_8 => UNWINDOWED_466 ,
										MUX_10_1_IN_9 => UNWINDOWED_466 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_233
									);
MUX_REORD_UNIT_234 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_234 ,
										MUX_10_1_IN_1 => UNWINDOWED_233 ,
										MUX_10_1_IN_2 => UNWINDOWED_236 ,
										MUX_10_1_IN_3 => UNWINDOWED_229 ,
										MUX_10_1_IN_4 => UNWINDOWED_244 ,
										MUX_10_1_IN_5 => UNWINDOWED_213 ,
										MUX_10_1_IN_6 => UNWINDOWED_213 ,
										MUX_10_1_IN_7 => UNWINDOWED_213 ,
										MUX_10_1_IN_8 => UNWINDOWED_468 ,
										MUX_10_1_IN_9 => UNWINDOWED_468 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_234
									);
MUX_REORD_UNIT_235 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_235 ,
										MUX_10_1_IN_1 => UNWINDOWED_235 ,
										MUX_10_1_IN_2 => UNWINDOWED_238 ,
										MUX_10_1_IN_3 => UNWINDOWED_231 ,
										MUX_10_1_IN_4 => UNWINDOWED_246 ,
										MUX_10_1_IN_5 => UNWINDOWED_215 ,
										MUX_10_1_IN_6 => UNWINDOWED_215 ,
										MUX_10_1_IN_7 => UNWINDOWED_215 ,
										MUX_10_1_IN_8 => UNWINDOWED_470 ,
										MUX_10_1_IN_9 => UNWINDOWED_470 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_235
									);
MUX_REORD_UNIT_236 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_236 ,
										MUX_10_1_IN_1 => UNWINDOWED_236 ,
										MUX_10_1_IN_2 => UNWINDOWED_233 ,
										MUX_10_1_IN_3 => UNWINDOWED_233 ,
										MUX_10_1_IN_4 => UNWINDOWED_248 ,
										MUX_10_1_IN_5 => UNWINDOWED_217 ,
										MUX_10_1_IN_6 => UNWINDOWED_217 ,
										MUX_10_1_IN_7 => UNWINDOWED_217 ,
										MUX_10_1_IN_8 => UNWINDOWED_472 ,
										MUX_10_1_IN_9 => UNWINDOWED_472 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_236
									);
MUX_REORD_UNIT_237 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_237 ,
										MUX_10_1_IN_1 => UNWINDOWED_238 ,
										MUX_10_1_IN_2 => UNWINDOWED_235 ,
										MUX_10_1_IN_3 => UNWINDOWED_235 ,
										MUX_10_1_IN_4 => UNWINDOWED_250 ,
										MUX_10_1_IN_5 => UNWINDOWED_219 ,
										MUX_10_1_IN_6 => UNWINDOWED_219 ,
										MUX_10_1_IN_7 => UNWINDOWED_219 ,
										MUX_10_1_IN_8 => UNWINDOWED_474 ,
										MUX_10_1_IN_9 => UNWINDOWED_474 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_237
									);
MUX_REORD_UNIT_238 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_238 ,
										MUX_10_1_IN_1 => UNWINDOWED_237 ,
										MUX_10_1_IN_2 => UNWINDOWED_237 ,
										MUX_10_1_IN_3 => UNWINDOWED_237 ,
										MUX_10_1_IN_4 => UNWINDOWED_252 ,
										MUX_10_1_IN_5 => UNWINDOWED_221 ,
										MUX_10_1_IN_6 => UNWINDOWED_221 ,
										MUX_10_1_IN_7 => UNWINDOWED_221 ,
										MUX_10_1_IN_8 => UNWINDOWED_476 ,
										MUX_10_1_IN_9 => UNWINDOWED_476 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_238
									);
MUX_REORD_UNIT_239 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_239 ,
										MUX_10_1_IN_1 => UNWINDOWED_239 ,
										MUX_10_1_IN_2 => UNWINDOWED_239 ,
										MUX_10_1_IN_3 => UNWINDOWED_239 ,
										MUX_10_1_IN_4 => UNWINDOWED_254 ,
										MUX_10_1_IN_5 => UNWINDOWED_223 ,
										MUX_10_1_IN_6 => UNWINDOWED_223 ,
										MUX_10_1_IN_7 => UNWINDOWED_223 ,
										MUX_10_1_IN_8 => UNWINDOWED_478 ,
										MUX_10_1_IN_9 => UNWINDOWED_478 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_239
									);
MUX_REORD_UNIT_240 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_240 ,
										MUX_10_1_IN_1 => UNWINDOWED_240 ,
										MUX_10_1_IN_2 => UNWINDOWED_240 ,
										MUX_10_1_IN_3 => UNWINDOWED_240 ,
										MUX_10_1_IN_4 => UNWINDOWED_225 ,
										MUX_10_1_IN_5 => UNWINDOWED_225 ,
										MUX_10_1_IN_6 => UNWINDOWED_225 ,
										MUX_10_1_IN_7 => UNWINDOWED_225 ,
										MUX_10_1_IN_8 => UNWINDOWED_480 ,
										MUX_10_1_IN_9 => UNWINDOWED_480 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_240
									);
MUX_REORD_UNIT_241 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_241 ,
										MUX_10_1_IN_1 => UNWINDOWED_242 ,
										MUX_10_1_IN_2 => UNWINDOWED_242 ,
										MUX_10_1_IN_3 => UNWINDOWED_242 ,
										MUX_10_1_IN_4 => UNWINDOWED_227 ,
										MUX_10_1_IN_5 => UNWINDOWED_227 ,
										MUX_10_1_IN_6 => UNWINDOWED_227 ,
										MUX_10_1_IN_7 => UNWINDOWED_227 ,
										MUX_10_1_IN_8 => UNWINDOWED_482 ,
										MUX_10_1_IN_9 => UNWINDOWED_482 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_241
									);
MUX_REORD_UNIT_242 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_242 ,
										MUX_10_1_IN_1 => UNWINDOWED_241 ,
										MUX_10_1_IN_2 => UNWINDOWED_244 ,
										MUX_10_1_IN_3 => UNWINDOWED_244 ,
										MUX_10_1_IN_4 => UNWINDOWED_229 ,
										MUX_10_1_IN_5 => UNWINDOWED_229 ,
										MUX_10_1_IN_6 => UNWINDOWED_229 ,
										MUX_10_1_IN_7 => UNWINDOWED_229 ,
										MUX_10_1_IN_8 => UNWINDOWED_484 ,
										MUX_10_1_IN_9 => UNWINDOWED_484 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_242
									);
MUX_REORD_UNIT_243 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_243 ,
										MUX_10_1_IN_1 => UNWINDOWED_243 ,
										MUX_10_1_IN_2 => UNWINDOWED_246 ,
										MUX_10_1_IN_3 => UNWINDOWED_246 ,
										MUX_10_1_IN_4 => UNWINDOWED_231 ,
										MUX_10_1_IN_5 => UNWINDOWED_231 ,
										MUX_10_1_IN_6 => UNWINDOWED_231 ,
										MUX_10_1_IN_7 => UNWINDOWED_231 ,
										MUX_10_1_IN_8 => UNWINDOWED_486 ,
										MUX_10_1_IN_9 => UNWINDOWED_486 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_243
									);
MUX_REORD_UNIT_244 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_244 ,
										MUX_10_1_IN_1 => UNWINDOWED_244 ,
										MUX_10_1_IN_2 => UNWINDOWED_241 ,
										MUX_10_1_IN_3 => UNWINDOWED_248 ,
										MUX_10_1_IN_4 => UNWINDOWED_233 ,
										MUX_10_1_IN_5 => UNWINDOWED_233 ,
										MUX_10_1_IN_6 => UNWINDOWED_233 ,
										MUX_10_1_IN_7 => UNWINDOWED_233 ,
										MUX_10_1_IN_8 => UNWINDOWED_488 ,
										MUX_10_1_IN_9 => UNWINDOWED_488 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_244
									);
MUX_REORD_UNIT_245 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_245 ,
										MUX_10_1_IN_1 => UNWINDOWED_246 ,
										MUX_10_1_IN_2 => UNWINDOWED_243 ,
										MUX_10_1_IN_3 => UNWINDOWED_250 ,
										MUX_10_1_IN_4 => UNWINDOWED_235 ,
										MUX_10_1_IN_5 => UNWINDOWED_235 ,
										MUX_10_1_IN_6 => UNWINDOWED_235 ,
										MUX_10_1_IN_7 => UNWINDOWED_235 ,
										MUX_10_1_IN_8 => UNWINDOWED_490 ,
										MUX_10_1_IN_9 => UNWINDOWED_490 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_245
									);
MUX_REORD_UNIT_246 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_246 ,
										MUX_10_1_IN_1 => UNWINDOWED_245 ,
										MUX_10_1_IN_2 => UNWINDOWED_245 ,
										MUX_10_1_IN_3 => UNWINDOWED_252 ,
										MUX_10_1_IN_4 => UNWINDOWED_237 ,
										MUX_10_1_IN_5 => UNWINDOWED_237 ,
										MUX_10_1_IN_6 => UNWINDOWED_237 ,
										MUX_10_1_IN_7 => UNWINDOWED_237 ,
										MUX_10_1_IN_8 => UNWINDOWED_492 ,
										MUX_10_1_IN_9 => UNWINDOWED_492 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_246
									);
MUX_REORD_UNIT_247 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_247 ,
										MUX_10_1_IN_1 => UNWINDOWED_247 ,
										MUX_10_1_IN_2 => UNWINDOWED_247 ,
										MUX_10_1_IN_3 => UNWINDOWED_254 ,
										MUX_10_1_IN_4 => UNWINDOWED_239 ,
										MUX_10_1_IN_5 => UNWINDOWED_239 ,
										MUX_10_1_IN_6 => UNWINDOWED_239 ,
										MUX_10_1_IN_7 => UNWINDOWED_239 ,
										MUX_10_1_IN_8 => UNWINDOWED_494 ,
										MUX_10_1_IN_9 => UNWINDOWED_494 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_247
									);
MUX_REORD_UNIT_248 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_248 ,
										MUX_10_1_IN_1 => UNWINDOWED_248 ,
										MUX_10_1_IN_2 => UNWINDOWED_248 ,
										MUX_10_1_IN_3 => UNWINDOWED_241 ,
										MUX_10_1_IN_4 => UNWINDOWED_241 ,
										MUX_10_1_IN_5 => UNWINDOWED_241 ,
										MUX_10_1_IN_6 => UNWINDOWED_241 ,
										MUX_10_1_IN_7 => UNWINDOWED_241 ,
										MUX_10_1_IN_8 => UNWINDOWED_496 ,
										MUX_10_1_IN_9 => UNWINDOWED_496 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_248
									);
MUX_REORD_UNIT_249 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_249 ,
										MUX_10_1_IN_1 => UNWINDOWED_250 ,
										MUX_10_1_IN_2 => UNWINDOWED_250 ,
										MUX_10_1_IN_3 => UNWINDOWED_243 ,
										MUX_10_1_IN_4 => UNWINDOWED_243 ,
										MUX_10_1_IN_5 => UNWINDOWED_243 ,
										MUX_10_1_IN_6 => UNWINDOWED_243 ,
										MUX_10_1_IN_7 => UNWINDOWED_243 ,
										MUX_10_1_IN_8 => UNWINDOWED_498 ,
										MUX_10_1_IN_9 => UNWINDOWED_498 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_249
									);
MUX_REORD_UNIT_250 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_250 ,
										MUX_10_1_IN_1 => UNWINDOWED_249 ,
										MUX_10_1_IN_2 => UNWINDOWED_252 ,
										MUX_10_1_IN_3 => UNWINDOWED_245 ,
										MUX_10_1_IN_4 => UNWINDOWED_245 ,
										MUX_10_1_IN_5 => UNWINDOWED_245 ,
										MUX_10_1_IN_6 => UNWINDOWED_245 ,
										MUX_10_1_IN_7 => UNWINDOWED_245 ,
										MUX_10_1_IN_8 => UNWINDOWED_500 ,
										MUX_10_1_IN_9 => UNWINDOWED_500 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_250
									);
MUX_REORD_UNIT_251 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_251 ,
										MUX_10_1_IN_1 => UNWINDOWED_251 ,
										MUX_10_1_IN_2 => UNWINDOWED_254 ,
										MUX_10_1_IN_3 => UNWINDOWED_247 ,
										MUX_10_1_IN_4 => UNWINDOWED_247 ,
										MUX_10_1_IN_5 => UNWINDOWED_247 ,
										MUX_10_1_IN_6 => UNWINDOWED_247 ,
										MUX_10_1_IN_7 => UNWINDOWED_247 ,
										MUX_10_1_IN_8 => UNWINDOWED_502 ,
										MUX_10_1_IN_9 => UNWINDOWED_502 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_251
									);
MUX_REORD_UNIT_252 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_252 ,
										MUX_10_1_IN_1 => UNWINDOWED_252 ,
										MUX_10_1_IN_2 => UNWINDOWED_249 ,
										MUX_10_1_IN_3 => UNWINDOWED_249 ,
										MUX_10_1_IN_4 => UNWINDOWED_249 ,
										MUX_10_1_IN_5 => UNWINDOWED_249 ,
										MUX_10_1_IN_6 => UNWINDOWED_249 ,
										MUX_10_1_IN_7 => UNWINDOWED_249 ,
										MUX_10_1_IN_8 => UNWINDOWED_504 ,
										MUX_10_1_IN_9 => UNWINDOWED_504 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_252
									);
MUX_REORD_UNIT_253 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_253 ,
										MUX_10_1_IN_1 => UNWINDOWED_254 ,
										MUX_10_1_IN_2 => UNWINDOWED_251 ,
										MUX_10_1_IN_3 => UNWINDOWED_251 ,
										MUX_10_1_IN_4 => UNWINDOWED_251 ,
										MUX_10_1_IN_5 => UNWINDOWED_251 ,
										MUX_10_1_IN_6 => UNWINDOWED_251 ,
										MUX_10_1_IN_7 => UNWINDOWED_251 ,
										MUX_10_1_IN_8 => UNWINDOWED_506 ,
										MUX_10_1_IN_9 => UNWINDOWED_506 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_253
									);
MUX_REORD_UNIT_254 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_254 ,
										MUX_10_1_IN_1 => UNWINDOWED_253 ,
										MUX_10_1_IN_2 => UNWINDOWED_253 ,
										MUX_10_1_IN_3 => UNWINDOWED_253 ,
										MUX_10_1_IN_4 => UNWINDOWED_253 ,
										MUX_10_1_IN_5 => UNWINDOWED_253 ,
										MUX_10_1_IN_6 => UNWINDOWED_253 ,
										MUX_10_1_IN_7 => UNWINDOWED_253 ,
										MUX_10_1_IN_8 => UNWINDOWED_508 ,
										MUX_10_1_IN_9 => UNWINDOWED_508 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_254
									);
MUX_REORD_UNIT_255 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_255 ,
										MUX_10_1_IN_1 => UNWINDOWED_255 ,
										MUX_10_1_IN_2 => UNWINDOWED_255 ,
										MUX_10_1_IN_3 => UNWINDOWED_255 ,
										MUX_10_1_IN_4 => UNWINDOWED_255 ,
										MUX_10_1_IN_5 => UNWINDOWED_255 ,
										MUX_10_1_IN_6 => UNWINDOWED_255 ,
										MUX_10_1_IN_7 => UNWINDOWED_255 ,
										MUX_10_1_IN_8 => UNWINDOWED_510 ,
										MUX_10_1_IN_9 => UNWINDOWED_510 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_255
									);
MUX_REORD_UNIT_256 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_256 ,
										MUX_10_1_IN_1 => UNWINDOWED_256 ,
										MUX_10_1_IN_2 => UNWINDOWED_256 ,
										MUX_10_1_IN_3 => UNWINDOWED_256 ,
										MUX_10_1_IN_4 => UNWINDOWED_256 ,
										MUX_10_1_IN_5 => UNWINDOWED_256 ,
										MUX_10_1_IN_6 => UNWINDOWED_256 ,
										MUX_10_1_IN_7 => UNWINDOWED_256 ,
										MUX_10_1_IN_8 => UNWINDOWED_1 ,
										MUX_10_1_IN_9 => UNWINDOWED_512 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_256
									);
MUX_REORD_UNIT_257 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_257 ,
										MUX_10_1_IN_1 => UNWINDOWED_258 ,
										MUX_10_1_IN_2 => UNWINDOWED_258 ,
										MUX_10_1_IN_3 => UNWINDOWED_258 ,
										MUX_10_1_IN_4 => UNWINDOWED_258 ,
										MUX_10_1_IN_5 => UNWINDOWED_258 ,
										MUX_10_1_IN_6 => UNWINDOWED_258 ,
										MUX_10_1_IN_7 => UNWINDOWED_258 ,
										MUX_10_1_IN_8 => UNWINDOWED_3 ,
										MUX_10_1_IN_9 => UNWINDOWED_514 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_257
									);
MUX_REORD_UNIT_258 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_258 ,
										MUX_10_1_IN_1 => UNWINDOWED_257 ,
										MUX_10_1_IN_2 => UNWINDOWED_260 ,
										MUX_10_1_IN_3 => UNWINDOWED_260 ,
										MUX_10_1_IN_4 => UNWINDOWED_260 ,
										MUX_10_1_IN_5 => UNWINDOWED_260 ,
										MUX_10_1_IN_6 => UNWINDOWED_260 ,
										MUX_10_1_IN_7 => UNWINDOWED_260 ,
										MUX_10_1_IN_8 => UNWINDOWED_5 ,
										MUX_10_1_IN_9 => UNWINDOWED_516 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_258
									);
MUX_REORD_UNIT_259 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_259 ,
										MUX_10_1_IN_1 => UNWINDOWED_259 ,
										MUX_10_1_IN_2 => UNWINDOWED_262 ,
										MUX_10_1_IN_3 => UNWINDOWED_262 ,
										MUX_10_1_IN_4 => UNWINDOWED_262 ,
										MUX_10_1_IN_5 => UNWINDOWED_262 ,
										MUX_10_1_IN_6 => UNWINDOWED_262 ,
										MUX_10_1_IN_7 => UNWINDOWED_262 ,
										MUX_10_1_IN_8 => UNWINDOWED_7 ,
										MUX_10_1_IN_9 => UNWINDOWED_518 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_259
									);
MUX_REORD_UNIT_260 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_260 ,
										MUX_10_1_IN_1 => UNWINDOWED_260 ,
										MUX_10_1_IN_2 => UNWINDOWED_257 ,
										MUX_10_1_IN_3 => UNWINDOWED_264 ,
										MUX_10_1_IN_4 => UNWINDOWED_264 ,
										MUX_10_1_IN_5 => UNWINDOWED_264 ,
										MUX_10_1_IN_6 => UNWINDOWED_264 ,
										MUX_10_1_IN_7 => UNWINDOWED_264 ,
										MUX_10_1_IN_8 => UNWINDOWED_9 ,
										MUX_10_1_IN_9 => UNWINDOWED_520 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_260
									);
MUX_REORD_UNIT_261 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_261 ,
										MUX_10_1_IN_1 => UNWINDOWED_262 ,
										MUX_10_1_IN_2 => UNWINDOWED_259 ,
										MUX_10_1_IN_3 => UNWINDOWED_266 ,
										MUX_10_1_IN_4 => UNWINDOWED_266 ,
										MUX_10_1_IN_5 => UNWINDOWED_266 ,
										MUX_10_1_IN_6 => UNWINDOWED_266 ,
										MUX_10_1_IN_7 => UNWINDOWED_266 ,
										MUX_10_1_IN_8 => UNWINDOWED_11 ,
										MUX_10_1_IN_9 => UNWINDOWED_522 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_261
									);
MUX_REORD_UNIT_262 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_262 ,
										MUX_10_1_IN_1 => UNWINDOWED_261 ,
										MUX_10_1_IN_2 => UNWINDOWED_261 ,
										MUX_10_1_IN_3 => UNWINDOWED_268 ,
										MUX_10_1_IN_4 => UNWINDOWED_268 ,
										MUX_10_1_IN_5 => UNWINDOWED_268 ,
										MUX_10_1_IN_6 => UNWINDOWED_268 ,
										MUX_10_1_IN_7 => UNWINDOWED_268 ,
										MUX_10_1_IN_8 => UNWINDOWED_13 ,
										MUX_10_1_IN_9 => UNWINDOWED_524 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_262
									);
MUX_REORD_UNIT_263 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_263 ,
										MUX_10_1_IN_1 => UNWINDOWED_263 ,
										MUX_10_1_IN_2 => UNWINDOWED_263 ,
										MUX_10_1_IN_3 => UNWINDOWED_270 ,
										MUX_10_1_IN_4 => UNWINDOWED_270 ,
										MUX_10_1_IN_5 => UNWINDOWED_270 ,
										MUX_10_1_IN_6 => UNWINDOWED_270 ,
										MUX_10_1_IN_7 => UNWINDOWED_270 ,
										MUX_10_1_IN_8 => UNWINDOWED_15 ,
										MUX_10_1_IN_9 => UNWINDOWED_526 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_263
									);
MUX_REORD_UNIT_264 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_264 ,
										MUX_10_1_IN_1 => UNWINDOWED_264 ,
										MUX_10_1_IN_2 => UNWINDOWED_264 ,
										MUX_10_1_IN_3 => UNWINDOWED_257 ,
										MUX_10_1_IN_4 => UNWINDOWED_272 ,
										MUX_10_1_IN_5 => UNWINDOWED_272 ,
										MUX_10_1_IN_6 => UNWINDOWED_272 ,
										MUX_10_1_IN_7 => UNWINDOWED_272 ,
										MUX_10_1_IN_8 => UNWINDOWED_17 ,
										MUX_10_1_IN_9 => UNWINDOWED_528 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_264
									);
MUX_REORD_UNIT_265 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_265 ,
										MUX_10_1_IN_1 => UNWINDOWED_266 ,
										MUX_10_1_IN_2 => UNWINDOWED_266 ,
										MUX_10_1_IN_3 => UNWINDOWED_259 ,
										MUX_10_1_IN_4 => UNWINDOWED_274 ,
										MUX_10_1_IN_5 => UNWINDOWED_274 ,
										MUX_10_1_IN_6 => UNWINDOWED_274 ,
										MUX_10_1_IN_7 => UNWINDOWED_274 ,
										MUX_10_1_IN_8 => UNWINDOWED_19 ,
										MUX_10_1_IN_9 => UNWINDOWED_530 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_265
									);
MUX_REORD_UNIT_266 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_266 ,
										MUX_10_1_IN_1 => UNWINDOWED_265 ,
										MUX_10_1_IN_2 => UNWINDOWED_268 ,
										MUX_10_1_IN_3 => UNWINDOWED_261 ,
										MUX_10_1_IN_4 => UNWINDOWED_276 ,
										MUX_10_1_IN_5 => UNWINDOWED_276 ,
										MUX_10_1_IN_6 => UNWINDOWED_276 ,
										MUX_10_1_IN_7 => UNWINDOWED_276 ,
										MUX_10_1_IN_8 => UNWINDOWED_21 ,
										MUX_10_1_IN_9 => UNWINDOWED_532 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_266
									);
MUX_REORD_UNIT_267 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_267 ,
										MUX_10_1_IN_1 => UNWINDOWED_267 ,
										MUX_10_1_IN_2 => UNWINDOWED_270 ,
										MUX_10_1_IN_3 => UNWINDOWED_263 ,
										MUX_10_1_IN_4 => UNWINDOWED_278 ,
										MUX_10_1_IN_5 => UNWINDOWED_278 ,
										MUX_10_1_IN_6 => UNWINDOWED_278 ,
										MUX_10_1_IN_7 => UNWINDOWED_278 ,
										MUX_10_1_IN_8 => UNWINDOWED_23 ,
										MUX_10_1_IN_9 => UNWINDOWED_534 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_267
									);
MUX_REORD_UNIT_268 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_268 ,
										MUX_10_1_IN_1 => UNWINDOWED_268 ,
										MUX_10_1_IN_2 => UNWINDOWED_265 ,
										MUX_10_1_IN_3 => UNWINDOWED_265 ,
										MUX_10_1_IN_4 => UNWINDOWED_280 ,
										MUX_10_1_IN_5 => UNWINDOWED_280 ,
										MUX_10_1_IN_6 => UNWINDOWED_280 ,
										MUX_10_1_IN_7 => UNWINDOWED_280 ,
										MUX_10_1_IN_8 => UNWINDOWED_25 ,
										MUX_10_1_IN_9 => UNWINDOWED_536 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_268
									);
MUX_REORD_UNIT_269 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_269 ,
										MUX_10_1_IN_1 => UNWINDOWED_270 ,
										MUX_10_1_IN_2 => UNWINDOWED_267 ,
										MUX_10_1_IN_3 => UNWINDOWED_267 ,
										MUX_10_1_IN_4 => UNWINDOWED_282 ,
										MUX_10_1_IN_5 => UNWINDOWED_282 ,
										MUX_10_1_IN_6 => UNWINDOWED_282 ,
										MUX_10_1_IN_7 => UNWINDOWED_282 ,
										MUX_10_1_IN_8 => UNWINDOWED_27 ,
										MUX_10_1_IN_9 => UNWINDOWED_538 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_269
									);
MUX_REORD_UNIT_270 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_270 ,
										MUX_10_1_IN_1 => UNWINDOWED_269 ,
										MUX_10_1_IN_2 => UNWINDOWED_269 ,
										MUX_10_1_IN_3 => UNWINDOWED_269 ,
										MUX_10_1_IN_4 => UNWINDOWED_284 ,
										MUX_10_1_IN_5 => UNWINDOWED_284 ,
										MUX_10_1_IN_6 => UNWINDOWED_284 ,
										MUX_10_1_IN_7 => UNWINDOWED_284 ,
										MUX_10_1_IN_8 => UNWINDOWED_29 ,
										MUX_10_1_IN_9 => UNWINDOWED_540 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_270
									);
MUX_REORD_UNIT_271 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_271 ,
										MUX_10_1_IN_1 => UNWINDOWED_271 ,
										MUX_10_1_IN_2 => UNWINDOWED_271 ,
										MUX_10_1_IN_3 => UNWINDOWED_271 ,
										MUX_10_1_IN_4 => UNWINDOWED_286 ,
										MUX_10_1_IN_5 => UNWINDOWED_286 ,
										MUX_10_1_IN_6 => UNWINDOWED_286 ,
										MUX_10_1_IN_7 => UNWINDOWED_286 ,
										MUX_10_1_IN_8 => UNWINDOWED_31 ,
										MUX_10_1_IN_9 => UNWINDOWED_542 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_271
									);
MUX_REORD_UNIT_272 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_272 ,
										MUX_10_1_IN_1 => UNWINDOWED_272 ,
										MUX_10_1_IN_2 => UNWINDOWED_272 ,
										MUX_10_1_IN_3 => UNWINDOWED_272 ,
										MUX_10_1_IN_4 => UNWINDOWED_257 ,
										MUX_10_1_IN_5 => UNWINDOWED_288 ,
										MUX_10_1_IN_6 => UNWINDOWED_288 ,
										MUX_10_1_IN_7 => UNWINDOWED_288 ,
										MUX_10_1_IN_8 => UNWINDOWED_33 ,
										MUX_10_1_IN_9 => UNWINDOWED_544 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_272
									);
MUX_REORD_UNIT_273 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_273 ,
										MUX_10_1_IN_1 => UNWINDOWED_274 ,
										MUX_10_1_IN_2 => UNWINDOWED_274 ,
										MUX_10_1_IN_3 => UNWINDOWED_274 ,
										MUX_10_1_IN_4 => UNWINDOWED_259 ,
										MUX_10_1_IN_5 => UNWINDOWED_290 ,
										MUX_10_1_IN_6 => UNWINDOWED_290 ,
										MUX_10_1_IN_7 => UNWINDOWED_290 ,
										MUX_10_1_IN_8 => UNWINDOWED_35 ,
										MUX_10_1_IN_9 => UNWINDOWED_546 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_273
									);
MUX_REORD_UNIT_274 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_274 ,
										MUX_10_1_IN_1 => UNWINDOWED_273 ,
										MUX_10_1_IN_2 => UNWINDOWED_276 ,
										MUX_10_1_IN_3 => UNWINDOWED_276 ,
										MUX_10_1_IN_4 => UNWINDOWED_261 ,
										MUX_10_1_IN_5 => UNWINDOWED_292 ,
										MUX_10_1_IN_6 => UNWINDOWED_292 ,
										MUX_10_1_IN_7 => UNWINDOWED_292 ,
										MUX_10_1_IN_8 => UNWINDOWED_37 ,
										MUX_10_1_IN_9 => UNWINDOWED_548 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_274
									);
MUX_REORD_UNIT_275 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_275 ,
										MUX_10_1_IN_1 => UNWINDOWED_275 ,
										MUX_10_1_IN_2 => UNWINDOWED_278 ,
										MUX_10_1_IN_3 => UNWINDOWED_278 ,
										MUX_10_1_IN_4 => UNWINDOWED_263 ,
										MUX_10_1_IN_5 => UNWINDOWED_294 ,
										MUX_10_1_IN_6 => UNWINDOWED_294 ,
										MUX_10_1_IN_7 => UNWINDOWED_294 ,
										MUX_10_1_IN_8 => UNWINDOWED_39 ,
										MUX_10_1_IN_9 => UNWINDOWED_550 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_275
									);
MUX_REORD_UNIT_276 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_276 ,
										MUX_10_1_IN_1 => UNWINDOWED_276 ,
										MUX_10_1_IN_2 => UNWINDOWED_273 ,
										MUX_10_1_IN_3 => UNWINDOWED_280 ,
										MUX_10_1_IN_4 => UNWINDOWED_265 ,
										MUX_10_1_IN_5 => UNWINDOWED_296 ,
										MUX_10_1_IN_6 => UNWINDOWED_296 ,
										MUX_10_1_IN_7 => UNWINDOWED_296 ,
										MUX_10_1_IN_8 => UNWINDOWED_41 ,
										MUX_10_1_IN_9 => UNWINDOWED_552 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_276
									);
MUX_REORD_UNIT_277 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_277 ,
										MUX_10_1_IN_1 => UNWINDOWED_278 ,
										MUX_10_1_IN_2 => UNWINDOWED_275 ,
										MUX_10_1_IN_3 => UNWINDOWED_282 ,
										MUX_10_1_IN_4 => UNWINDOWED_267 ,
										MUX_10_1_IN_5 => UNWINDOWED_298 ,
										MUX_10_1_IN_6 => UNWINDOWED_298 ,
										MUX_10_1_IN_7 => UNWINDOWED_298 ,
										MUX_10_1_IN_8 => UNWINDOWED_43 ,
										MUX_10_1_IN_9 => UNWINDOWED_554 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_277
									);
MUX_REORD_UNIT_278 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_278 ,
										MUX_10_1_IN_1 => UNWINDOWED_277 ,
										MUX_10_1_IN_2 => UNWINDOWED_277 ,
										MUX_10_1_IN_3 => UNWINDOWED_284 ,
										MUX_10_1_IN_4 => UNWINDOWED_269 ,
										MUX_10_1_IN_5 => UNWINDOWED_300 ,
										MUX_10_1_IN_6 => UNWINDOWED_300 ,
										MUX_10_1_IN_7 => UNWINDOWED_300 ,
										MUX_10_1_IN_8 => UNWINDOWED_45 ,
										MUX_10_1_IN_9 => UNWINDOWED_556 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_278
									);
MUX_REORD_UNIT_279 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_279 ,
										MUX_10_1_IN_1 => UNWINDOWED_279 ,
										MUX_10_1_IN_2 => UNWINDOWED_279 ,
										MUX_10_1_IN_3 => UNWINDOWED_286 ,
										MUX_10_1_IN_4 => UNWINDOWED_271 ,
										MUX_10_1_IN_5 => UNWINDOWED_302 ,
										MUX_10_1_IN_6 => UNWINDOWED_302 ,
										MUX_10_1_IN_7 => UNWINDOWED_302 ,
										MUX_10_1_IN_8 => UNWINDOWED_47 ,
										MUX_10_1_IN_9 => UNWINDOWED_558 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_279
									);
MUX_REORD_UNIT_280 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_280 ,
										MUX_10_1_IN_1 => UNWINDOWED_280 ,
										MUX_10_1_IN_2 => UNWINDOWED_280 ,
										MUX_10_1_IN_3 => UNWINDOWED_273 ,
										MUX_10_1_IN_4 => UNWINDOWED_273 ,
										MUX_10_1_IN_5 => UNWINDOWED_304 ,
										MUX_10_1_IN_6 => UNWINDOWED_304 ,
										MUX_10_1_IN_7 => UNWINDOWED_304 ,
										MUX_10_1_IN_8 => UNWINDOWED_49 ,
										MUX_10_1_IN_9 => UNWINDOWED_560 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_280
									);
MUX_REORD_UNIT_281 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_281 ,
										MUX_10_1_IN_1 => UNWINDOWED_282 ,
										MUX_10_1_IN_2 => UNWINDOWED_282 ,
										MUX_10_1_IN_3 => UNWINDOWED_275 ,
										MUX_10_1_IN_4 => UNWINDOWED_275 ,
										MUX_10_1_IN_5 => UNWINDOWED_306 ,
										MUX_10_1_IN_6 => UNWINDOWED_306 ,
										MUX_10_1_IN_7 => UNWINDOWED_306 ,
										MUX_10_1_IN_8 => UNWINDOWED_51 ,
										MUX_10_1_IN_9 => UNWINDOWED_562 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_281
									);
MUX_REORD_UNIT_282 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_282 ,
										MUX_10_1_IN_1 => UNWINDOWED_281 ,
										MUX_10_1_IN_2 => UNWINDOWED_284 ,
										MUX_10_1_IN_3 => UNWINDOWED_277 ,
										MUX_10_1_IN_4 => UNWINDOWED_277 ,
										MUX_10_1_IN_5 => UNWINDOWED_308 ,
										MUX_10_1_IN_6 => UNWINDOWED_308 ,
										MUX_10_1_IN_7 => UNWINDOWED_308 ,
										MUX_10_1_IN_8 => UNWINDOWED_53 ,
										MUX_10_1_IN_9 => UNWINDOWED_564 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_282
									);
MUX_REORD_UNIT_283 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_283 ,
										MUX_10_1_IN_1 => UNWINDOWED_283 ,
										MUX_10_1_IN_2 => UNWINDOWED_286 ,
										MUX_10_1_IN_3 => UNWINDOWED_279 ,
										MUX_10_1_IN_4 => UNWINDOWED_279 ,
										MUX_10_1_IN_5 => UNWINDOWED_310 ,
										MUX_10_1_IN_6 => UNWINDOWED_310 ,
										MUX_10_1_IN_7 => UNWINDOWED_310 ,
										MUX_10_1_IN_8 => UNWINDOWED_55 ,
										MUX_10_1_IN_9 => UNWINDOWED_566 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_283
									);
MUX_REORD_UNIT_284 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_284 ,
										MUX_10_1_IN_1 => UNWINDOWED_284 ,
										MUX_10_1_IN_2 => UNWINDOWED_281 ,
										MUX_10_1_IN_3 => UNWINDOWED_281 ,
										MUX_10_1_IN_4 => UNWINDOWED_281 ,
										MUX_10_1_IN_5 => UNWINDOWED_312 ,
										MUX_10_1_IN_6 => UNWINDOWED_312 ,
										MUX_10_1_IN_7 => UNWINDOWED_312 ,
										MUX_10_1_IN_8 => UNWINDOWED_57 ,
										MUX_10_1_IN_9 => UNWINDOWED_568 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_284
									);
MUX_REORD_UNIT_285 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_285 ,
										MUX_10_1_IN_1 => UNWINDOWED_286 ,
										MUX_10_1_IN_2 => UNWINDOWED_283 ,
										MUX_10_1_IN_3 => UNWINDOWED_283 ,
										MUX_10_1_IN_4 => UNWINDOWED_283 ,
										MUX_10_1_IN_5 => UNWINDOWED_314 ,
										MUX_10_1_IN_6 => UNWINDOWED_314 ,
										MUX_10_1_IN_7 => UNWINDOWED_314 ,
										MUX_10_1_IN_8 => UNWINDOWED_59 ,
										MUX_10_1_IN_9 => UNWINDOWED_570 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_285
									);
MUX_REORD_UNIT_286 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_286 ,
										MUX_10_1_IN_1 => UNWINDOWED_285 ,
										MUX_10_1_IN_2 => UNWINDOWED_285 ,
										MUX_10_1_IN_3 => UNWINDOWED_285 ,
										MUX_10_1_IN_4 => UNWINDOWED_285 ,
										MUX_10_1_IN_5 => UNWINDOWED_316 ,
										MUX_10_1_IN_6 => UNWINDOWED_316 ,
										MUX_10_1_IN_7 => UNWINDOWED_316 ,
										MUX_10_1_IN_8 => UNWINDOWED_61 ,
										MUX_10_1_IN_9 => UNWINDOWED_572 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_286
									);
MUX_REORD_UNIT_287 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_287 ,
										MUX_10_1_IN_1 => UNWINDOWED_287 ,
										MUX_10_1_IN_2 => UNWINDOWED_287 ,
										MUX_10_1_IN_3 => UNWINDOWED_287 ,
										MUX_10_1_IN_4 => UNWINDOWED_287 ,
										MUX_10_1_IN_5 => UNWINDOWED_318 ,
										MUX_10_1_IN_6 => UNWINDOWED_318 ,
										MUX_10_1_IN_7 => UNWINDOWED_318 ,
										MUX_10_1_IN_8 => UNWINDOWED_63 ,
										MUX_10_1_IN_9 => UNWINDOWED_574 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_287
									);
MUX_REORD_UNIT_288 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_288 ,
										MUX_10_1_IN_1 => UNWINDOWED_288 ,
										MUX_10_1_IN_2 => UNWINDOWED_288 ,
										MUX_10_1_IN_3 => UNWINDOWED_288 ,
										MUX_10_1_IN_4 => UNWINDOWED_288 ,
										MUX_10_1_IN_5 => UNWINDOWED_257 ,
										MUX_10_1_IN_6 => UNWINDOWED_320 ,
										MUX_10_1_IN_7 => UNWINDOWED_320 ,
										MUX_10_1_IN_8 => UNWINDOWED_65 ,
										MUX_10_1_IN_9 => UNWINDOWED_576 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_288
									);
MUX_REORD_UNIT_289 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_289 ,
										MUX_10_1_IN_1 => UNWINDOWED_290 ,
										MUX_10_1_IN_2 => UNWINDOWED_290 ,
										MUX_10_1_IN_3 => UNWINDOWED_290 ,
										MUX_10_1_IN_4 => UNWINDOWED_290 ,
										MUX_10_1_IN_5 => UNWINDOWED_259 ,
										MUX_10_1_IN_6 => UNWINDOWED_322 ,
										MUX_10_1_IN_7 => UNWINDOWED_322 ,
										MUX_10_1_IN_8 => UNWINDOWED_67 ,
										MUX_10_1_IN_9 => UNWINDOWED_578 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_289
									);
MUX_REORD_UNIT_290 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_290 ,
										MUX_10_1_IN_1 => UNWINDOWED_289 ,
										MUX_10_1_IN_2 => UNWINDOWED_292 ,
										MUX_10_1_IN_3 => UNWINDOWED_292 ,
										MUX_10_1_IN_4 => UNWINDOWED_292 ,
										MUX_10_1_IN_5 => UNWINDOWED_261 ,
										MUX_10_1_IN_6 => UNWINDOWED_324 ,
										MUX_10_1_IN_7 => UNWINDOWED_324 ,
										MUX_10_1_IN_8 => UNWINDOWED_69 ,
										MUX_10_1_IN_9 => UNWINDOWED_580 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_290
									);
MUX_REORD_UNIT_291 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_291 ,
										MUX_10_1_IN_1 => UNWINDOWED_291 ,
										MUX_10_1_IN_2 => UNWINDOWED_294 ,
										MUX_10_1_IN_3 => UNWINDOWED_294 ,
										MUX_10_1_IN_4 => UNWINDOWED_294 ,
										MUX_10_1_IN_5 => UNWINDOWED_263 ,
										MUX_10_1_IN_6 => UNWINDOWED_326 ,
										MUX_10_1_IN_7 => UNWINDOWED_326 ,
										MUX_10_1_IN_8 => UNWINDOWED_71 ,
										MUX_10_1_IN_9 => UNWINDOWED_582 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_291
									);
MUX_REORD_UNIT_292 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_292 ,
										MUX_10_1_IN_1 => UNWINDOWED_292 ,
										MUX_10_1_IN_2 => UNWINDOWED_289 ,
										MUX_10_1_IN_3 => UNWINDOWED_296 ,
										MUX_10_1_IN_4 => UNWINDOWED_296 ,
										MUX_10_1_IN_5 => UNWINDOWED_265 ,
										MUX_10_1_IN_6 => UNWINDOWED_328 ,
										MUX_10_1_IN_7 => UNWINDOWED_328 ,
										MUX_10_1_IN_8 => UNWINDOWED_73 ,
										MUX_10_1_IN_9 => UNWINDOWED_584 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_292
									);
MUX_REORD_UNIT_293 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_293 ,
										MUX_10_1_IN_1 => UNWINDOWED_294 ,
										MUX_10_1_IN_2 => UNWINDOWED_291 ,
										MUX_10_1_IN_3 => UNWINDOWED_298 ,
										MUX_10_1_IN_4 => UNWINDOWED_298 ,
										MUX_10_1_IN_5 => UNWINDOWED_267 ,
										MUX_10_1_IN_6 => UNWINDOWED_330 ,
										MUX_10_1_IN_7 => UNWINDOWED_330 ,
										MUX_10_1_IN_8 => UNWINDOWED_75 ,
										MUX_10_1_IN_9 => UNWINDOWED_586 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_293
									);
MUX_REORD_UNIT_294 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_294 ,
										MUX_10_1_IN_1 => UNWINDOWED_293 ,
										MUX_10_1_IN_2 => UNWINDOWED_293 ,
										MUX_10_1_IN_3 => UNWINDOWED_300 ,
										MUX_10_1_IN_4 => UNWINDOWED_300 ,
										MUX_10_1_IN_5 => UNWINDOWED_269 ,
										MUX_10_1_IN_6 => UNWINDOWED_332 ,
										MUX_10_1_IN_7 => UNWINDOWED_332 ,
										MUX_10_1_IN_8 => UNWINDOWED_77 ,
										MUX_10_1_IN_9 => UNWINDOWED_588 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_294
									);
MUX_REORD_UNIT_295 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_295 ,
										MUX_10_1_IN_1 => UNWINDOWED_295 ,
										MUX_10_1_IN_2 => UNWINDOWED_295 ,
										MUX_10_1_IN_3 => UNWINDOWED_302 ,
										MUX_10_1_IN_4 => UNWINDOWED_302 ,
										MUX_10_1_IN_5 => UNWINDOWED_271 ,
										MUX_10_1_IN_6 => UNWINDOWED_334 ,
										MUX_10_1_IN_7 => UNWINDOWED_334 ,
										MUX_10_1_IN_8 => UNWINDOWED_79 ,
										MUX_10_1_IN_9 => UNWINDOWED_590 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_295
									);
MUX_REORD_UNIT_296 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_296 ,
										MUX_10_1_IN_1 => UNWINDOWED_296 ,
										MUX_10_1_IN_2 => UNWINDOWED_296 ,
										MUX_10_1_IN_3 => UNWINDOWED_289 ,
										MUX_10_1_IN_4 => UNWINDOWED_304 ,
										MUX_10_1_IN_5 => UNWINDOWED_273 ,
										MUX_10_1_IN_6 => UNWINDOWED_336 ,
										MUX_10_1_IN_7 => UNWINDOWED_336 ,
										MUX_10_1_IN_8 => UNWINDOWED_81 ,
										MUX_10_1_IN_9 => UNWINDOWED_592 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_296
									);
MUX_REORD_UNIT_297 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_297 ,
										MUX_10_1_IN_1 => UNWINDOWED_298 ,
										MUX_10_1_IN_2 => UNWINDOWED_298 ,
										MUX_10_1_IN_3 => UNWINDOWED_291 ,
										MUX_10_1_IN_4 => UNWINDOWED_306 ,
										MUX_10_1_IN_5 => UNWINDOWED_275 ,
										MUX_10_1_IN_6 => UNWINDOWED_338 ,
										MUX_10_1_IN_7 => UNWINDOWED_338 ,
										MUX_10_1_IN_8 => UNWINDOWED_83 ,
										MUX_10_1_IN_9 => UNWINDOWED_594 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_297
									);
MUX_REORD_UNIT_298 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_298 ,
										MUX_10_1_IN_1 => UNWINDOWED_297 ,
										MUX_10_1_IN_2 => UNWINDOWED_300 ,
										MUX_10_1_IN_3 => UNWINDOWED_293 ,
										MUX_10_1_IN_4 => UNWINDOWED_308 ,
										MUX_10_1_IN_5 => UNWINDOWED_277 ,
										MUX_10_1_IN_6 => UNWINDOWED_340 ,
										MUX_10_1_IN_7 => UNWINDOWED_340 ,
										MUX_10_1_IN_8 => UNWINDOWED_85 ,
										MUX_10_1_IN_9 => UNWINDOWED_596 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_298
									);
MUX_REORD_UNIT_299 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_299 ,
										MUX_10_1_IN_1 => UNWINDOWED_299 ,
										MUX_10_1_IN_2 => UNWINDOWED_302 ,
										MUX_10_1_IN_3 => UNWINDOWED_295 ,
										MUX_10_1_IN_4 => UNWINDOWED_310 ,
										MUX_10_1_IN_5 => UNWINDOWED_279 ,
										MUX_10_1_IN_6 => UNWINDOWED_342 ,
										MUX_10_1_IN_7 => UNWINDOWED_342 ,
										MUX_10_1_IN_8 => UNWINDOWED_87 ,
										MUX_10_1_IN_9 => UNWINDOWED_598 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_299
									);
MUX_REORD_UNIT_300 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_300 ,
										MUX_10_1_IN_1 => UNWINDOWED_300 ,
										MUX_10_1_IN_2 => UNWINDOWED_297 ,
										MUX_10_1_IN_3 => UNWINDOWED_297 ,
										MUX_10_1_IN_4 => UNWINDOWED_312 ,
										MUX_10_1_IN_5 => UNWINDOWED_281 ,
										MUX_10_1_IN_6 => UNWINDOWED_344 ,
										MUX_10_1_IN_7 => UNWINDOWED_344 ,
										MUX_10_1_IN_8 => UNWINDOWED_89 ,
										MUX_10_1_IN_9 => UNWINDOWED_600 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_300
									);
MUX_REORD_UNIT_301 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_301 ,
										MUX_10_1_IN_1 => UNWINDOWED_302 ,
										MUX_10_1_IN_2 => UNWINDOWED_299 ,
										MUX_10_1_IN_3 => UNWINDOWED_299 ,
										MUX_10_1_IN_4 => UNWINDOWED_314 ,
										MUX_10_1_IN_5 => UNWINDOWED_283 ,
										MUX_10_1_IN_6 => UNWINDOWED_346 ,
										MUX_10_1_IN_7 => UNWINDOWED_346 ,
										MUX_10_1_IN_8 => UNWINDOWED_91 ,
										MUX_10_1_IN_9 => UNWINDOWED_602 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_301
									);
MUX_REORD_UNIT_302 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_302 ,
										MUX_10_1_IN_1 => UNWINDOWED_301 ,
										MUX_10_1_IN_2 => UNWINDOWED_301 ,
										MUX_10_1_IN_3 => UNWINDOWED_301 ,
										MUX_10_1_IN_4 => UNWINDOWED_316 ,
										MUX_10_1_IN_5 => UNWINDOWED_285 ,
										MUX_10_1_IN_6 => UNWINDOWED_348 ,
										MUX_10_1_IN_7 => UNWINDOWED_348 ,
										MUX_10_1_IN_8 => UNWINDOWED_93 ,
										MUX_10_1_IN_9 => UNWINDOWED_604 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_302
									);
MUX_REORD_UNIT_303 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_303 ,
										MUX_10_1_IN_1 => UNWINDOWED_303 ,
										MUX_10_1_IN_2 => UNWINDOWED_303 ,
										MUX_10_1_IN_3 => UNWINDOWED_303 ,
										MUX_10_1_IN_4 => UNWINDOWED_318 ,
										MUX_10_1_IN_5 => UNWINDOWED_287 ,
										MUX_10_1_IN_6 => UNWINDOWED_350 ,
										MUX_10_1_IN_7 => UNWINDOWED_350 ,
										MUX_10_1_IN_8 => UNWINDOWED_95 ,
										MUX_10_1_IN_9 => UNWINDOWED_606 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_303
									);
MUX_REORD_UNIT_304 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_304 ,
										MUX_10_1_IN_1 => UNWINDOWED_304 ,
										MUX_10_1_IN_2 => UNWINDOWED_304 ,
										MUX_10_1_IN_3 => UNWINDOWED_304 ,
										MUX_10_1_IN_4 => UNWINDOWED_289 ,
										MUX_10_1_IN_5 => UNWINDOWED_289 ,
										MUX_10_1_IN_6 => UNWINDOWED_352 ,
										MUX_10_1_IN_7 => UNWINDOWED_352 ,
										MUX_10_1_IN_8 => UNWINDOWED_97 ,
										MUX_10_1_IN_9 => UNWINDOWED_608 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_304
									);
MUX_REORD_UNIT_305 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_305 ,
										MUX_10_1_IN_1 => UNWINDOWED_306 ,
										MUX_10_1_IN_2 => UNWINDOWED_306 ,
										MUX_10_1_IN_3 => UNWINDOWED_306 ,
										MUX_10_1_IN_4 => UNWINDOWED_291 ,
										MUX_10_1_IN_5 => UNWINDOWED_291 ,
										MUX_10_1_IN_6 => UNWINDOWED_354 ,
										MUX_10_1_IN_7 => UNWINDOWED_354 ,
										MUX_10_1_IN_8 => UNWINDOWED_99 ,
										MUX_10_1_IN_9 => UNWINDOWED_610 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_305
									);
MUX_REORD_UNIT_306 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_306 ,
										MUX_10_1_IN_1 => UNWINDOWED_305 ,
										MUX_10_1_IN_2 => UNWINDOWED_308 ,
										MUX_10_1_IN_3 => UNWINDOWED_308 ,
										MUX_10_1_IN_4 => UNWINDOWED_293 ,
										MUX_10_1_IN_5 => UNWINDOWED_293 ,
										MUX_10_1_IN_6 => UNWINDOWED_356 ,
										MUX_10_1_IN_7 => UNWINDOWED_356 ,
										MUX_10_1_IN_8 => UNWINDOWED_101 ,
										MUX_10_1_IN_9 => UNWINDOWED_612 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_306
									);
MUX_REORD_UNIT_307 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_307 ,
										MUX_10_1_IN_1 => UNWINDOWED_307 ,
										MUX_10_1_IN_2 => UNWINDOWED_310 ,
										MUX_10_1_IN_3 => UNWINDOWED_310 ,
										MUX_10_1_IN_4 => UNWINDOWED_295 ,
										MUX_10_1_IN_5 => UNWINDOWED_295 ,
										MUX_10_1_IN_6 => UNWINDOWED_358 ,
										MUX_10_1_IN_7 => UNWINDOWED_358 ,
										MUX_10_1_IN_8 => UNWINDOWED_103 ,
										MUX_10_1_IN_9 => UNWINDOWED_614 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_307
									);
MUX_REORD_UNIT_308 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_308 ,
										MUX_10_1_IN_1 => UNWINDOWED_308 ,
										MUX_10_1_IN_2 => UNWINDOWED_305 ,
										MUX_10_1_IN_3 => UNWINDOWED_312 ,
										MUX_10_1_IN_4 => UNWINDOWED_297 ,
										MUX_10_1_IN_5 => UNWINDOWED_297 ,
										MUX_10_1_IN_6 => UNWINDOWED_360 ,
										MUX_10_1_IN_7 => UNWINDOWED_360 ,
										MUX_10_1_IN_8 => UNWINDOWED_105 ,
										MUX_10_1_IN_9 => UNWINDOWED_616 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_308
									);
MUX_REORD_UNIT_309 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_309 ,
										MUX_10_1_IN_1 => UNWINDOWED_310 ,
										MUX_10_1_IN_2 => UNWINDOWED_307 ,
										MUX_10_1_IN_3 => UNWINDOWED_314 ,
										MUX_10_1_IN_4 => UNWINDOWED_299 ,
										MUX_10_1_IN_5 => UNWINDOWED_299 ,
										MUX_10_1_IN_6 => UNWINDOWED_362 ,
										MUX_10_1_IN_7 => UNWINDOWED_362 ,
										MUX_10_1_IN_8 => UNWINDOWED_107 ,
										MUX_10_1_IN_9 => UNWINDOWED_618 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_309
									);
MUX_REORD_UNIT_310 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_310 ,
										MUX_10_1_IN_1 => UNWINDOWED_309 ,
										MUX_10_1_IN_2 => UNWINDOWED_309 ,
										MUX_10_1_IN_3 => UNWINDOWED_316 ,
										MUX_10_1_IN_4 => UNWINDOWED_301 ,
										MUX_10_1_IN_5 => UNWINDOWED_301 ,
										MUX_10_1_IN_6 => UNWINDOWED_364 ,
										MUX_10_1_IN_7 => UNWINDOWED_364 ,
										MUX_10_1_IN_8 => UNWINDOWED_109 ,
										MUX_10_1_IN_9 => UNWINDOWED_620 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_310
									);
MUX_REORD_UNIT_311 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_311 ,
										MUX_10_1_IN_1 => UNWINDOWED_311 ,
										MUX_10_1_IN_2 => UNWINDOWED_311 ,
										MUX_10_1_IN_3 => UNWINDOWED_318 ,
										MUX_10_1_IN_4 => UNWINDOWED_303 ,
										MUX_10_1_IN_5 => UNWINDOWED_303 ,
										MUX_10_1_IN_6 => UNWINDOWED_366 ,
										MUX_10_1_IN_7 => UNWINDOWED_366 ,
										MUX_10_1_IN_8 => UNWINDOWED_111 ,
										MUX_10_1_IN_9 => UNWINDOWED_622 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_311
									);
MUX_REORD_UNIT_312 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_312 ,
										MUX_10_1_IN_1 => UNWINDOWED_312 ,
										MUX_10_1_IN_2 => UNWINDOWED_312 ,
										MUX_10_1_IN_3 => UNWINDOWED_305 ,
										MUX_10_1_IN_4 => UNWINDOWED_305 ,
										MUX_10_1_IN_5 => UNWINDOWED_305 ,
										MUX_10_1_IN_6 => UNWINDOWED_368 ,
										MUX_10_1_IN_7 => UNWINDOWED_368 ,
										MUX_10_1_IN_8 => UNWINDOWED_113 ,
										MUX_10_1_IN_9 => UNWINDOWED_624 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_312
									);
MUX_REORD_UNIT_313 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_313 ,
										MUX_10_1_IN_1 => UNWINDOWED_314 ,
										MUX_10_1_IN_2 => UNWINDOWED_314 ,
										MUX_10_1_IN_3 => UNWINDOWED_307 ,
										MUX_10_1_IN_4 => UNWINDOWED_307 ,
										MUX_10_1_IN_5 => UNWINDOWED_307 ,
										MUX_10_1_IN_6 => UNWINDOWED_370 ,
										MUX_10_1_IN_7 => UNWINDOWED_370 ,
										MUX_10_1_IN_8 => UNWINDOWED_115 ,
										MUX_10_1_IN_9 => UNWINDOWED_626 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_313
									);
MUX_REORD_UNIT_314 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_314 ,
										MUX_10_1_IN_1 => UNWINDOWED_313 ,
										MUX_10_1_IN_2 => UNWINDOWED_316 ,
										MUX_10_1_IN_3 => UNWINDOWED_309 ,
										MUX_10_1_IN_4 => UNWINDOWED_309 ,
										MUX_10_1_IN_5 => UNWINDOWED_309 ,
										MUX_10_1_IN_6 => UNWINDOWED_372 ,
										MUX_10_1_IN_7 => UNWINDOWED_372 ,
										MUX_10_1_IN_8 => UNWINDOWED_117 ,
										MUX_10_1_IN_9 => UNWINDOWED_628 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_314
									);
MUX_REORD_UNIT_315 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_315 ,
										MUX_10_1_IN_1 => UNWINDOWED_315 ,
										MUX_10_1_IN_2 => UNWINDOWED_318 ,
										MUX_10_1_IN_3 => UNWINDOWED_311 ,
										MUX_10_1_IN_4 => UNWINDOWED_311 ,
										MUX_10_1_IN_5 => UNWINDOWED_311 ,
										MUX_10_1_IN_6 => UNWINDOWED_374 ,
										MUX_10_1_IN_7 => UNWINDOWED_374 ,
										MUX_10_1_IN_8 => UNWINDOWED_119 ,
										MUX_10_1_IN_9 => UNWINDOWED_630 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_315
									);
MUX_REORD_UNIT_316 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_316 ,
										MUX_10_1_IN_1 => UNWINDOWED_316 ,
										MUX_10_1_IN_2 => UNWINDOWED_313 ,
										MUX_10_1_IN_3 => UNWINDOWED_313 ,
										MUX_10_1_IN_4 => UNWINDOWED_313 ,
										MUX_10_1_IN_5 => UNWINDOWED_313 ,
										MUX_10_1_IN_6 => UNWINDOWED_376 ,
										MUX_10_1_IN_7 => UNWINDOWED_376 ,
										MUX_10_1_IN_8 => UNWINDOWED_121 ,
										MUX_10_1_IN_9 => UNWINDOWED_632 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_316
									);
MUX_REORD_UNIT_317 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_317 ,
										MUX_10_1_IN_1 => UNWINDOWED_318 ,
										MUX_10_1_IN_2 => UNWINDOWED_315 ,
										MUX_10_1_IN_3 => UNWINDOWED_315 ,
										MUX_10_1_IN_4 => UNWINDOWED_315 ,
										MUX_10_1_IN_5 => UNWINDOWED_315 ,
										MUX_10_1_IN_6 => UNWINDOWED_378 ,
										MUX_10_1_IN_7 => UNWINDOWED_378 ,
										MUX_10_1_IN_8 => UNWINDOWED_123 ,
										MUX_10_1_IN_9 => UNWINDOWED_634 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_317
									);
MUX_REORD_UNIT_318 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_318 ,
										MUX_10_1_IN_1 => UNWINDOWED_317 ,
										MUX_10_1_IN_2 => UNWINDOWED_317 ,
										MUX_10_1_IN_3 => UNWINDOWED_317 ,
										MUX_10_1_IN_4 => UNWINDOWED_317 ,
										MUX_10_1_IN_5 => UNWINDOWED_317 ,
										MUX_10_1_IN_6 => UNWINDOWED_380 ,
										MUX_10_1_IN_7 => UNWINDOWED_380 ,
										MUX_10_1_IN_8 => UNWINDOWED_125 ,
										MUX_10_1_IN_9 => UNWINDOWED_636 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_318
									);
MUX_REORD_UNIT_319 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_319 ,
										MUX_10_1_IN_1 => UNWINDOWED_319 ,
										MUX_10_1_IN_2 => UNWINDOWED_319 ,
										MUX_10_1_IN_3 => UNWINDOWED_319 ,
										MUX_10_1_IN_4 => UNWINDOWED_319 ,
										MUX_10_1_IN_5 => UNWINDOWED_319 ,
										MUX_10_1_IN_6 => UNWINDOWED_382 ,
										MUX_10_1_IN_7 => UNWINDOWED_382 ,
										MUX_10_1_IN_8 => UNWINDOWED_127 ,
										MUX_10_1_IN_9 => UNWINDOWED_638 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_319
									);
MUX_REORD_UNIT_320 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_320 ,
										MUX_10_1_IN_1 => UNWINDOWED_320 ,
										MUX_10_1_IN_2 => UNWINDOWED_320 ,
										MUX_10_1_IN_3 => UNWINDOWED_320 ,
										MUX_10_1_IN_4 => UNWINDOWED_320 ,
										MUX_10_1_IN_5 => UNWINDOWED_320 ,
										MUX_10_1_IN_6 => UNWINDOWED_257 ,
										MUX_10_1_IN_7 => UNWINDOWED_384 ,
										MUX_10_1_IN_8 => UNWINDOWED_129 ,
										MUX_10_1_IN_9 => UNWINDOWED_640 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_320
									);
MUX_REORD_UNIT_321 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_321 ,
										MUX_10_1_IN_1 => UNWINDOWED_322 ,
										MUX_10_1_IN_2 => UNWINDOWED_322 ,
										MUX_10_1_IN_3 => UNWINDOWED_322 ,
										MUX_10_1_IN_4 => UNWINDOWED_322 ,
										MUX_10_1_IN_5 => UNWINDOWED_322 ,
										MUX_10_1_IN_6 => UNWINDOWED_259 ,
										MUX_10_1_IN_7 => UNWINDOWED_386 ,
										MUX_10_1_IN_8 => UNWINDOWED_131 ,
										MUX_10_1_IN_9 => UNWINDOWED_642 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_321
									);
MUX_REORD_UNIT_322 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_322 ,
										MUX_10_1_IN_1 => UNWINDOWED_321 ,
										MUX_10_1_IN_2 => UNWINDOWED_324 ,
										MUX_10_1_IN_3 => UNWINDOWED_324 ,
										MUX_10_1_IN_4 => UNWINDOWED_324 ,
										MUX_10_1_IN_5 => UNWINDOWED_324 ,
										MUX_10_1_IN_6 => UNWINDOWED_261 ,
										MUX_10_1_IN_7 => UNWINDOWED_388 ,
										MUX_10_1_IN_8 => UNWINDOWED_133 ,
										MUX_10_1_IN_9 => UNWINDOWED_644 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_322
									);
MUX_REORD_UNIT_323 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_323 ,
										MUX_10_1_IN_1 => UNWINDOWED_323 ,
										MUX_10_1_IN_2 => UNWINDOWED_326 ,
										MUX_10_1_IN_3 => UNWINDOWED_326 ,
										MUX_10_1_IN_4 => UNWINDOWED_326 ,
										MUX_10_1_IN_5 => UNWINDOWED_326 ,
										MUX_10_1_IN_6 => UNWINDOWED_263 ,
										MUX_10_1_IN_7 => UNWINDOWED_390 ,
										MUX_10_1_IN_8 => UNWINDOWED_135 ,
										MUX_10_1_IN_9 => UNWINDOWED_646 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_323
									);
MUX_REORD_UNIT_324 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_324 ,
										MUX_10_1_IN_1 => UNWINDOWED_324 ,
										MUX_10_1_IN_2 => UNWINDOWED_321 ,
										MUX_10_1_IN_3 => UNWINDOWED_328 ,
										MUX_10_1_IN_4 => UNWINDOWED_328 ,
										MUX_10_1_IN_5 => UNWINDOWED_328 ,
										MUX_10_1_IN_6 => UNWINDOWED_265 ,
										MUX_10_1_IN_7 => UNWINDOWED_392 ,
										MUX_10_1_IN_8 => UNWINDOWED_137 ,
										MUX_10_1_IN_9 => UNWINDOWED_648 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_324
									);
MUX_REORD_UNIT_325 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_325 ,
										MUX_10_1_IN_1 => UNWINDOWED_326 ,
										MUX_10_1_IN_2 => UNWINDOWED_323 ,
										MUX_10_1_IN_3 => UNWINDOWED_330 ,
										MUX_10_1_IN_4 => UNWINDOWED_330 ,
										MUX_10_1_IN_5 => UNWINDOWED_330 ,
										MUX_10_1_IN_6 => UNWINDOWED_267 ,
										MUX_10_1_IN_7 => UNWINDOWED_394 ,
										MUX_10_1_IN_8 => UNWINDOWED_139 ,
										MUX_10_1_IN_9 => UNWINDOWED_650 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_325
									);
MUX_REORD_UNIT_326 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_326 ,
										MUX_10_1_IN_1 => UNWINDOWED_325 ,
										MUX_10_1_IN_2 => UNWINDOWED_325 ,
										MUX_10_1_IN_3 => UNWINDOWED_332 ,
										MUX_10_1_IN_4 => UNWINDOWED_332 ,
										MUX_10_1_IN_5 => UNWINDOWED_332 ,
										MUX_10_1_IN_6 => UNWINDOWED_269 ,
										MUX_10_1_IN_7 => UNWINDOWED_396 ,
										MUX_10_1_IN_8 => UNWINDOWED_141 ,
										MUX_10_1_IN_9 => UNWINDOWED_652 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_326
									);
MUX_REORD_UNIT_327 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_327 ,
										MUX_10_1_IN_1 => UNWINDOWED_327 ,
										MUX_10_1_IN_2 => UNWINDOWED_327 ,
										MUX_10_1_IN_3 => UNWINDOWED_334 ,
										MUX_10_1_IN_4 => UNWINDOWED_334 ,
										MUX_10_1_IN_5 => UNWINDOWED_334 ,
										MUX_10_1_IN_6 => UNWINDOWED_271 ,
										MUX_10_1_IN_7 => UNWINDOWED_398 ,
										MUX_10_1_IN_8 => UNWINDOWED_143 ,
										MUX_10_1_IN_9 => UNWINDOWED_654 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_327
									);
MUX_REORD_UNIT_328 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_328 ,
										MUX_10_1_IN_1 => UNWINDOWED_328 ,
										MUX_10_1_IN_2 => UNWINDOWED_328 ,
										MUX_10_1_IN_3 => UNWINDOWED_321 ,
										MUX_10_1_IN_4 => UNWINDOWED_336 ,
										MUX_10_1_IN_5 => UNWINDOWED_336 ,
										MUX_10_1_IN_6 => UNWINDOWED_273 ,
										MUX_10_1_IN_7 => UNWINDOWED_400 ,
										MUX_10_1_IN_8 => UNWINDOWED_145 ,
										MUX_10_1_IN_9 => UNWINDOWED_656 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_328
									);
MUX_REORD_UNIT_329 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_329 ,
										MUX_10_1_IN_1 => UNWINDOWED_330 ,
										MUX_10_1_IN_2 => UNWINDOWED_330 ,
										MUX_10_1_IN_3 => UNWINDOWED_323 ,
										MUX_10_1_IN_4 => UNWINDOWED_338 ,
										MUX_10_1_IN_5 => UNWINDOWED_338 ,
										MUX_10_1_IN_6 => UNWINDOWED_275 ,
										MUX_10_1_IN_7 => UNWINDOWED_402 ,
										MUX_10_1_IN_8 => UNWINDOWED_147 ,
										MUX_10_1_IN_9 => UNWINDOWED_658 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_329
									);
MUX_REORD_UNIT_330 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_330 ,
										MUX_10_1_IN_1 => UNWINDOWED_329 ,
										MUX_10_1_IN_2 => UNWINDOWED_332 ,
										MUX_10_1_IN_3 => UNWINDOWED_325 ,
										MUX_10_1_IN_4 => UNWINDOWED_340 ,
										MUX_10_1_IN_5 => UNWINDOWED_340 ,
										MUX_10_1_IN_6 => UNWINDOWED_277 ,
										MUX_10_1_IN_7 => UNWINDOWED_404 ,
										MUX_10_1_IN_8 => UNWINDOWED_149 ,
										MUX_10_1_IN_9 => UNWINDOWED_660 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_330
									);
MUX_REORD_UNIT_331 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_331 ,
										MUX_10_1_IN_1 => UNWINDOWED_331 ,
										MUX_10_1_IN_2 => UNWINDOWED_334 ,
										MUX_10_1_IN_3 => UNWINDOWED_327 ,
										MUX_10_1_IN_4 => UNWINDOWED_342 ,
										MUX_10_1_IN_5 => UNWINDOWED_342 ,
										MUX_10_1_IN_6 => UNWINDOWED_279 ,
										MUX_10_1_IN_7 => UNWINDOWED_406 ,
										MUX_10_1_IN_8 => UNWINDOWED_151 ,
										MUX_10_1_IN_9 => UNWINDOWED_662 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_331
									);
MUX_REORD_UNIT_332 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_332 ,
										MUX_10_1_IN_1 => UNWINDOWED_332 ,
										MUX_10_1_IN_2 => UNWINDOWED_329 ,
										MUX_10_1_IN_3 => UNWINDOWED_329 ,
										MUX_10_1_IN_4 => UNWINDOWED_344 ,
										MUX_10_1_IN_5 => UNWINDOWED_344 ,
										MUX_10_1_IN_6 => UNWINDOWED_281 ,
										MUX_10_1_IN_7 => UNWINDOWED_408 ,
										MUX_10_1_IN_8 => UNWINDOWED_153 ,
										MUX_10_1_IN_9 => UNWINDOWED_664 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_332
									);
MUX_REORD_UNIT_333 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_333 ,
										MUX_10_1_IN_1 => UNWINDOWED_334 ,
										MUX_10_1_IN_2 => UNWINDOWED_331 ,
										MUX_10_1_IN_3 => UNWINDOWED_331 ,
										MUX_10_1_IN_4 => UNWINDOWED_346 ,
										MUX_10_1_IN_5 => UNWINDOWED_346 ,
										MUX_10_1_IN_6 => UNWINDOWED_283 ,
										MUX_10_1_IN_7 => UNWINDOWED_410 ,
										MUX_10_1_IN_8 => UNWINDOWED_155 ,
										MUX_10_1_IN_9 => UNWINDOWED_666 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_333
									);
MUX_REORD_UNIT_334 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_334 ,
										MUX_10_1_IN_1 => UNWINDOWED_333 ,
										MUX_10_1_IN_2 => UNWINDOWED_333 ,
										MUX_10_1_IN_3 => UNWINDOWED_333 ,
										MUX_10_1_IN_4 => UNWINDOWED_348 ,
										MUX_10_1_IN_5 => UNWINDOWED_348 ,
										MUX_10_1_IN_6 => UNWINDOWED_285 ,
										MUX_10_1_IN_7 => UNWINDOWED_412 ,
										MUX_10_1_IN_8 => UNWINDOWED_157 ,
										MUX_10_1_IN_9 => UNWINDOWED_668 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_334
									);
MUX_REORD_UNIT_335 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_335 ,
										MUX_10_1_IN_1 => UNWINDOWED_335 ,
										MUX_10_1_IN_2 => UNWINDOWED_335 ,
										MUX_10_1_IN_3 => UNWINDOWED_335 ,
										MUX_10_1_IN_4 => UNWINDOWED_350 ,
										MUX_10_1_IN_5 => UNWINDOWED_350 ,
										MUX_10_1_IN_6 => UNWINDOWED_287 ,
										MUX_10_1_IN_7 => UNWINDOWED_414 ,
										MUX_10_1_IN_8 => UNWINDOWED_159 ,
										MUX_10_1_IN_9 => UNWINDOWED_670 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_335
									);
MUX_REORD_UNIT_336 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_336 ,
										MUX_10_1_IN_1 => UNWINDOWED_336 ,
										MUX_10_1_IN_2 => UNWINDOWED_336 ,
										MUX_10_1_IN_3 => UNWINDOWED_336 ,
										MUX_10_1_IN_4 => UNWINDOWED_321 ,
										MUX_10_1_IN_5 => UNWINDOWED_352 ,
										MUX_10_1_IN_6 => UNWINDOWED_289 ,
										MUX_10_1_IN_7 => UNWINDOWED_416 ,
										MUX_10_1_IN_8 => UNWINDOWED_161 ,
										MUX_10_1_IN_9 => UNWINDOWED_672 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_336
									);
MUX_REORD_UNIT_337 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_337 ,
										MUX_10_1_IN_1 => UNWINDOWED_338 ,
										MUX_10_1_IN_2 => UNWINDOWED_338 ,
										MUX_10_1_IN_3 => UNWINDOWED_338 ,
										MUX_10_1_IN_4 => UNWINDOWED_323 ,
										MUX_10_1_IN_5 => UNWINDOWED_354 ,
										MUX_10_1_IN_6 => UNWINDOWED_291 ,
										MUX_10_1_IN_7 => UNWINDOWED_418 ,
										MUX_10_1_IN_8 => UNWINDOWED_163 ,
										MUX_10_1_IN_9 => UNWINDOWED_674 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_337
									);
MUX_REORD_UNIT_338 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_338 ,
										MUX_10_1_IN_1 => UNWINDOWED_337 ,
										MUX_10_1_IN_2 => UNWINDOWED_340 ,
										MUX_10_1_IN_3 => UNWINDOWED_340 ,
										MUX_10_1_IN_4 => UNWINDOWED_325 ,
										MUX_10_1_IN_5 => UNWINDOWED_356 ,
										MUX_10_1_IN_6 => UNWINDOWED_293 ,
										MUX_10_1_IN_7 => UNWINDOWED_420 ,
										MUX_10_1_IN_8 => UNWINDOWED_165 ,
										MUX_10_1_IN_9 => UNWINDOWED_676 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_338
									);
MUX_REORD_UNIT_339 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_339 ,
										MUX_10_1_IN_1 => UNWINDOWED_339 ,
										MUX_10_1_IN_2 => UNWINDOWED_342 ,
										MUX_10_1_IN_3 => UNWINDOWED_342 ,
										MUX_10_1_IN_4 => UNWINDOWED_327 ,
										MUX_10_1_IN_5 => UNWINDOWED_358 ,
										MUX_10_1_IN_6 => UNWINDOWED_295 ,
										MUX_10_1_IN_7 => UNWINDOWED_422 ,
										MUX_10_1_IN_8 => UNWINDOWED_167 ,
										MUX_10_1_IN_9 => UNWINDOWED_678 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_339
									);
MUX_REORD_UNIT_340 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_340 ,
										MUX_10_1_IN_1 => UNWINDOWED_340 ,
										MUX_10_1_IN_2 => UNWINDOWED_337 ,
										MUX_10_1_IN_3 => UNWINDOWED_344 ,
										MUX_10_1_IN_4 => UNWINDOWED_329 ,
										MUX_10_1_IN_5 => UNWINDOWED_360 ,
										MUX_10_1_IN_6 => UNWINDOWED_297 ,
										MUX_10_1_IN_7 => UNWINDOWED_424 ,
										MUX_10_1_IN_8 => UNWINDOWED_169 ,
										MUX_10_1_IN_9 => UNWINDOWED_680 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_340
									);
MUX_REORD_UNIT_341 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_341 ,
										MUX_10_1_IN_1 => UNWINDOWED_342 ,
										MUX_10_1_IN_2 => UNWINDOWED_339 ,
										MUX_10_1_IN_3 => UNWINDOWED_346 ,
										MUX_10_1_IN_4 => UNWINDOWED_331 ,
										MUX_10_1_IN_5 => UNWINDOWED_362 ,
										MUX_10_1_IN_6 => UNWINDOWED_299 ,
										MUX_10_1_IN_7 => UNWINDOWED_426 ,
										MUX_10_1_IN_8 => UNWINDOWED_171 ,
										MUX_10_1_IN_9 => UNWINDOWED_682 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_341
									);
MUX_REORD_UNIT_342 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_342 ,
										MUX_10_1_IN_1 => UNWINDOWED_341 ,
										MUX_10_1_IN_2 => UNWINDOWED_341 ,
										MUX_10_1_IN_3 => UNWINDOWED_348 ,
										MUX_10_1_IN_4 => UNWINDOWED_333 ,
										MUX_10_1_IN_5 => UNWINDOWED_364 ,
										MUX_10_1_IN_6 => UNWINDOWED_301 ,
										MUX_10_1_IN_7 => UNWINDOWED_428 ,
										MUX_10_1_IN_8 => UNWINDOWED_173 ,
										MUX_10_1_IN_9 => UNWINDOWED_684 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_342
									);
MUX_REORD_UNIT_343 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_343 ,
										MUX_10_1_IN_1 => UNWINDOWED_343 ,
										MUX_10_1_IN_2 => UNWINDOWED_343 ,
										MUX_10_1_IN_3 => UNWINDOWED_350 ,
										MUX_10_1_IN_4 => UNWINDOWED_335 ,
										MUX_10_1_IN_5 => UNWINDOWED_366 ,
										MUX_10_1_IN_6 => UNWINDOWED_303 ,
										MUX_10_1_IN_7 => UNWINDOWED_430 ,
										MUX_10_1_IN_8 => UNWINDOWED_175 ,
										MUX_10_1_IN_9 => UNWINDOWED_686 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_343
									);
MUX_REORD_UNIT_344 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_344 ,
										MUX_10_1_IN_1 => UNWINDOWED_344 ,
										MUX_10_1_IN_2 => UNWINDOWED_344 ,
										MUX_10_1_IN_3 => UNWINDOWED_337 ,
										MUX_10_1_IN_4 => UNWINDOWED_337 ,
										MUX_10_1_IN_5 => UNWINDOWED_368 ,
										MUX_10_1_IN_6 => UNWINDOWED_305 ,
										MUX_10_1_IN_7 => UNWINDOWED_432 ,
										MUX_10_1_IN_8 => UNWINDOWED_177 ,
										MUX_10_1_IN_9 => UNWINDOWED_688 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_344
									);
MUX_REORD_UNIT_345 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_345 ,
										MUX_10_1_IN_1 => UNWINDOWED_346 ,
										MUX_10_1_IN_2 => UNWINDOWED_346 ,
										MUX_10_1_IN_3 => UNWINDOWED_339 ,
										MUX_10_1_IN_4 => UNWINDOWED_339 ,
										MUX_10_1_IN_5 => UNWINDOWED_370 ,
										MUX_10_1_IN_6 => UNWINDOWED_307 ,
										MUX_10_1_IN_7 => UNWINDOWED_434 ,
										MUX_10_1_IN_8 => UNWINDOWED_179 ,
										MUX_10_1_IN_9 => UNWINDOWED_690 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_345
									);
MUX_REORD_UNIT_346 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_346 ,
										MUX_10_1_IN_1 => UNWINDOWED_345 ,
										MUX_10_1_IN_2 => UNWINDOWED_348 ,
										MUX_10_1_IN_3 => UNWINDOWED_341 ,
										MUX_10_1_IN_4 => UNWINDOWED_341 ,
										MUX_10_1_IN_5 => UNWINDOWED_372 ,
										MUX_10_1_IN_6 => UNWINDOWED_309 ,
										MUX_10_1_IN_7 => UNWINDOWED_436 ,
										MUX_10_1_IN_8 => UNWINDOWED_181 ,
										MUX_10_1_IN_9 => UNWINDOWED_692 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_346
									);
MUX_REORD_UNIT_347 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_347 ,
										MUX_10_1_IN_1 => UNWINDOWED_347 ,
										MUX_10_1_IN_2 => UNWINDOWED_350 ,
										MUX_10_1_IN_3 => UNWINDOWED_343 ,
										MUX_10_1_IN_4 => UNWINDOWED_343 ,
										MUX_10_1_IN_5 => UNWINDOWED_374 ,
										MUX_10_1_IN_6 => UNWINDOWED_311 ,
										MUX_10_1_IN_7 => UNWINDOWED_438 ,
										MUX_10_1_IN_8 => UNWINDOWED_183 ,
										MUX_10_1_IN_9 => UNWINDOWED_694 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_347
									);
MUX_REORD_UNIT_348 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_348 ,
										MUX_10_1_IN_1 => UNWINDOWED_348 ,
										MUX_10_1_IN_2 => UNWINDOWED_345 ,
										MUX_10_1_IN_3 => UNWINDOWED_345 ,
										MUX_10_1_IN_4 => UNWINDOWED_345 ,
										MUX_10_1_IN_5 => UNWINDOWED_376 ,
										MUX_10_1_IN_6 => UNWINDOWED_313 ,
										MUX_10_1_IN_7 => UNWINDOWED_440 ,
										MUX_10_1_IN_8 => UNWINDOWED_185 ,
										MUX_10_1_IN_9 => UNWINDOWED_696 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_348
									);
MUX_REORD_UNIT_349 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_349 ,
										MUX_10_1_IN_1 => UNWINDOWED_350 ,
										MUX_10_1_IN_2 => UNWINDOWED_347 ,
										MUX_10_1_IN_3 => UNWINDOWED_347 ,
										MUX_10_1_IN_4 => UNWINDOWED_347 ,
										MUX_10_1_IN_5 => UNWINDOWED_378 ,
										MUX_10_1_IN_6 => UNWINDOWED_315 ,
										MUX_10_1_IN_7 => UNWINDOWED_442 ,
										MUX_10_1_IN_8 => UNWINDOWED_187 ,
										MUX_10_1_IN_9 => UNWINDOWED_698 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_349
									);
MUX_REORD_UNIT_350 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_350 ,
										MUX_10_1_IN_1 => UNWINDOWED_349 ,
										MUX_10_1_IN_2 => UNWINDOWED_349 ,
										MUX_10_1_IN_3 => UNWINDOWED_349 ,
										MUX_10_1_IN_4 => UNWINDOWED_349 ,
										MUX_10_1_IN_5 => UNWINDOWED_380 ,
										MUX_10_1_IN_6 => UNWINDOWED_317 ,
										MUX_10_1_IN_7 => UNWINDOWED_444 ,
										MUX_10_1_IN_8 => UNWINDOWED_189 ,
										MUX_10_1_IN_9 => UNWINDOWED_700 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_350
									);
MUX_REORD_UNIT_351 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_351 ,
										MUX_10_1_IN_1 => UNWINDOWED_351 ,
										MUX_10_1_IN_2 => UNWINDOWED_351 ,
										MUX_10_1_IN_3 => UNWINDOWED_351 ,
										MUX_10_1_IN_4 => UNWINDOWED_351 ,
										MUX_10_1_IN_5 => UNWINDOWED_382 ,
										MUX_10_1_IN_6 => UNWINDOWED_319 ,
										MUX_10_1_IN_7 => UNWINDOWED_446 ,
										MUX_10_1_IN_8 => UNWINDOWED_191 ,
										MUX_10_1_IN_9 => UNWINDOWED_702 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_351
									);
MUX_REORD_UNIT_352 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_352 ,
										MUX_10_1_IN_1 => UNWINDOWED_352 ,
										MUX_10_1_IN_2 => UNWINDOWED_352 ,
										MUX_10_1_IN_3 => UNWINDOWED_352 ,
										MUX_10_1_IN_4 => UNWINDOWED_352 ,
										MUX_10_1_IN_5 => UNWINDOWED_321 ,
										MUX_10_1_IN_6 => UNWINDOWED_321 ,
										MUX_10_1_IN_7 => UNWINDOWED_448 ,
										MUX_10_1_IN_8 => UNWINDOWED_193 ,
										MUX_10_1_IN_9 => UNWINDOWED_704 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_352
									);
MUX_REORD_UNIT_353 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_353 ,
										MUX_10_1_IN_1 => UNWINDOWED_354 ,
										MUX_10_1_IN_2 => UNWINDOWED_354 ,
										MUX_10_1_IN_3 => UNWINDOWED_354 ,
										MUX_10_1_IN_4 => UNWINDOWED_354 ,
										MUX_10_1_IN_5 => UNWINDOWED_323 ,
										MUX_10_1_IN_6 => UNWINDOWED_323 ,
										MUX_10_1_IN_7 => UNWINDOWED_450 ,
										MUX_10_1_IN_8 => UNWINDOWED_195 ,
										MUX_10_1_IN_9 => UNWINDOWED_706 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_353
									);
MUX_REORD_UNIT_354 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_354 ,
										MUX_10_1_IN_1 => UNWINDOWED_353 ,
										MUX_10_1_IN_2 => UNWINDOWED_356 ,
										MUX_10_1_IN_3 => UNWINDOWED_356 ,
										MUX_10_1_IN_4 => UNWINDOWED_356 ,
										MUX_10_1_IN_5 => UNWINDOWED_325 ,
										MUX_10_1_IN_6 => UNWINDOWED_325 ,
										MUX_10_1_IN_7 => UNWINDOWED_452 ,
										MUX_10_1_IN_8 => UNWINDOWED_197 ,
										MUX_10_1_IN_9 => UNWINDOWED_708 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_354
									);
MUX_REORD_UNIT_355 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_355 ,
										MUX_10_1_IN_1 => UNWINDOWED_355 ,
										MUX_10_1_IN_2 => UNWINDOWED_358 ,
										MUX_10_1_IN_3 => UNWINDOWED_358 ,
										MUX_10_1_IN_4 => UNWINDOWED_358 ,
										MUX_10_1_IN_5 => UNWINDOWED_327 ,
										MUX_10_1_IN_6 => UNWINDOWED_327 ,
										MUX_10_1_IN_7 => UNWINDOWED_454 ,
										MUX_10_1_IN_8 => UNWINDOWED_199 ,
										MUX_10_1_IN_9 => UNWINDOWED_710 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_355
									);
MUX_REORD_UNIT_356 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_356 ,
										MUX_10_1_IN_1 => UNWINDOWED_356 ,
										MUX_10_1_IN_2 => UNWINDOWED_353 ,
										MUX_10_1_IN_3 => UNWINDOWED_360 ,
										MUX_10_1_IN_4 => UNWINDOWED_360 ,
										MUX_10_1_IN_5 => UNWINDOWED_329 ,
										MUX_10_1_IN_6 => UNWINDOWED_329 ,
										MUX_10_1_IN_7 => UNWINDOWED_456 ,
										MUX_10_1_IN_8 => UNWINDOWED_201 ,
										MUX_10_1_IN_9 => UNWINDOWED_712 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_356
									);
MUX_REORD_UNIT_357 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_357 ,
										MUX_10_1_IN_1 => UNWINDOWED_358 ,
										MUX_10_1_IN_2 => UNWINDOWED_355 ,
										MUX_10_1_IN_3 => UNWINDOWED_362 ,
										MUX_10_1_IN_4 => UNWINDOWED_362 ,
										MUX_10_1_IN_5 => UNWINDOWED_331 ,
										MUX_10_1_IN_6 => UNWINDOWED_331 ,
										MUX_10_1_IN_7 => UNWINDOWED_458 ,
										MUX_10_1_IN_8 => UNWINDOWED_203 ,
										MUX_10_1_IN_9 => UNWINDOWED_714 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_357
									);
MUX_REORD_UNIT_358 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_358 ,
										MUX_10_1_IN_1 => UNWINDOWED_357 ,
										MUX_10_1_IN_2 => UNWINDOWED_357 ,
										MUX_10_1_IN_3 => UNWINDOWED_364 ,
										MUX_10_1_IN_4 => UNWINDOWED_364 ,
										MUX_10_1_IN_5 => UNWINDOWED_333 ,
										MUX_10_1_IN_6 => UNWINDOWED_333 ,
										MUX_10_1_IN_7 => UNWINDOWED_460 ,
										MUX_10_1_IN_8 => UNWINDOWED_205 ,
										MUX_10_1_IN_9 => UNWINDOWED_716 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_358
									);
MUX_REORD_UNIT_359 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_359 ,
										MUX_10_1_IN_1 => UNWINDOWED_359 ,
										MUX_10_1_IN_2 => UNWINDOWED_359 ,
										MUX_10_1_IN_3 => UNWINDOWED_366 ,
										MUX_10_1_IN_4 => UNWINDOWED_366 ,
										MUX_10_1_IN_5 => UNWINDOWED_335 ,
										MUX_10_1_IN_6 => UNWINDOWED_335 ,
										MUX_10_1_IN_7 => UNWINDOWED_462 ,
										MUX_10_1_IN_8 => UNWINDOWED_207 ,
										MUX_10_1_IN_9 => UNWINDOWED_718 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_359
									);
MUX_REORD_UNIT_360 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_360 ,
										MUX_10_1_IN_1 => UNWINDOWED_360 ,
										MUX_10_1_IN_2 => UNWINDOWED_360 ,
										MUX_10_1_IN_3 => UNWINDOWED_353 ,
										MUX_10_1_IN_4 => UNWINDOWED_368 ,
										MUX_10_1_IN_5 => UNWINDOWED_337 ,
										MUX_10_1_IN_6 => UNWINDOWED_337 ,
										MUX_10_1_IN_7 => UNWINDOWED_464 ,
										MUX_10_1_IN_8 => UNWINDOWED_209 ,
										MUX_10_1_IN_9 => UNWINDOWED_720 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_360
									);
MUX_REORD_UNIT_361 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_361 ,
										MUX_10_1_IN_1 => UNWINDOWED_362 ,
										MUX_10_1_IN_2 => UNWINDOWED_362 ,
										MUX_10_1_IN_3 => UNWINDOWED_355 ,
										MUX_10_1_IN_4 => UNWINDOWED_370 ,
										MUX_10_1_IN_5 => UNWINDOWED_339 ,
										MUX_10_1_IN_6 => UNWINDOWED_339 ,
										MUX_10_1_IN_7 => UNWINDOWED_466 ,
										MUX_10_1_IN_8 => UNWINDOWED_211 ,
										MUX_10_1_IN_9 => UNWINDOWED_722 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_361
									);
MUX_REORD_UNIT_362 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_362 ,
										MUX_10_1_IN_1 => UNWINDOWED_361 ,
										MUX_10_1_IN_2 => UNWINDOWED_364 ,
										MUX_10_1_IN_3 => UNWINDOWED_357 ,
										MUX_10_1_IN_4 => UNWINDOWED_372 ,
										MUX_10_1_IN_5 => UNWINDOWED_341 ,
										MUX_10_1_IN_6 => UNWINDOWED_341 ,
										MUX_10_1_IN_7 => UNWINDOWED_468 ,
										MUX_10_1_IN_8 => UNWINDOWED_213 ,
										MUX_10_1_IN_9 => UNWINDOWED_724 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_362
									);
MUX_REORD_UNIT_363 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_363 ,
										MUX_10_1_IN_1 => UNWINDOWED_363 ,
										MUX_10_1_IN_2 => UNWINDOWED_366 ,
										MUX_10_1_IN_3 => UNWINDOWED_359 ,
										MUX_10_1_IN_4 => UNWINDOWED_374 ,
										MUX_10_1_IN_5 => UNWINDOWED_343 ,
										MUX_10_1_IN_6 => UNWINDOWED_343 ,
										MUX_10_1_IN_7 => UNWINDOWED_470 ,
										MUX_10_1_IN_8 => UNWINDOWED_215 ,
										MUX_10_1_IN_9 => UNWINDOWED_726 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_363
									);
MUX_REORD_UNIT_364 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_364 ,
										MUX_10_1_IN_1 => UNWINDOWED_364 ,
										MUX_10_1_IN_2 => UNWINDOWED_361 ,
										MUX_10_1_IN_3 => UNWINDOWED_361 ,
										MUX_10_1_IN_4 => UNWINDOWED_376 ,
										MUX_10_1_IN_5 => UNWINDOWED_345 ,
										MUX_10_1_IN_6 => UNWINDOWED_345 ,
										MUX_10_1_IN_7 => UNWINDOWED_472 ,
										MUX_10_1_IN_8 => UNWINDOWED_217 ,
										MUX_10_1_IN_9 => UNWINDOWED_728 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_364
									);
MUX_REORD_UNIT_365 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_365 ,
										MUX_10_1_IN_1 => UNWINDOWED_366 ,
										MUX_10_1_IN_2 => UNWINDOWED_363 ,
										MUX_10_1_IN_3 => UNWINDOWED_363 ,
										MUX_10_1_IN_4 => UNWINDOWED_378 ,
										MUX_10_1_IN_5 => UNWINDOWED_347 ,
										MUX_10_1_IN_6 => UNWINDOWED_347 ,
										MUX_10_1_IN_7 => UNWINDOWED_474 ,
										MUX_10_1_IN_8 => UNWINDOWED_219 ,
										MUX_10_1_IN_9 => UNWINDOWED_730 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_365
									);
MUX_REORD_UNIT_366 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_366 ,
										MUX_10_1_IN_1 => UNWINDOWED_365 ,
										MUX_10_1_IN_2 => UNWINDOWED_365 ,
										MUX_10_1_IN_3 => UNWINDOWED_365 ,
										MUX_10_1_IN_4 => UNWINDOWED_380 ,
										MUX_10_1_IN_5 => UNWINDOWED_349 ,
										MUX_10_1_IN_6 => UNWINDOWED_349 ,
										MUX_10_1_IN_7 => UNWINDOWED_476 ,
										MUX_10_1_IN_8 => UNWINDOWED_221 ,
										MUX_10_1_IN_9 => UNWINDOWED_732 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_366
									);
MUX_REORD_UNIT_367 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_367 ,
										MUX_10_1_IN_1 => UNWINDOWED_367 ,
										MUX_10_1_IN_2 => UNWINDOWED_367 ,
										MUX_10_1_IN_3 => UNWINDOWED_367 ,
										MUX_10_1_IN_4 => UNWINDOWED_382 ,
										MUX_10_1_IN_5 => UNWINDOWED_351 ,
										MUX_10_1_IN_6 => UNWINDOWED_351 ,
										MUX_10_1_IN_7 => UNWINDOWED_478 ,
										MUX_10_1_IN_8 => UNWINDOWED_223 ,
										MUX_10_1_IN_9 => UNWINDOWED_734 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_367
									);
MUX_REORD_UNIT_368 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_368 ,
										MUX_10_1_IN_1 => UNWINDOWED_368 ,
										MUX_10_1_IN_2 => UNWINDOWED_368 ,
										MUX_10_1_IN_3 => UNWINDOWED_368 ,
										MUX_10_1_IN_4 => UNWINDOWED_353 ,
										MUX_10_1_IN_5 => UNWINDOWED_353 ,
										MUX_10_1_IN_6 => UNWINDOWED_353 ,
										MUX_10_1_IN_7 => UNWINDOWED_480 ,
										MUX_10_1_IN_8 => UNWINDOWED_225 ,
										MUX_10_1_IN_9 => UNWINDOWED_736 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_368
									);
MUX_REORD_UNIT_369 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_369 ,
										MUX_10_1_IN_1 => UNWINDOWED_370 ,
										MUX_10_1_IN_2 => UNWINDOWED_370 ,
										MUX_10_1_IN_3 => UNWINDOWED_370 ,
										MUX_10_1_IN_4 => UNWINDOWED_355 ,
										MUX_10_1_IN_5 => UNWINDOWED_355 ,
										MUX_10_1_IN_6 => UNWINDOWED_355 ,
										MUX_10_1_IN_7 => UNWINDOWED_482 ,
										MUX_10_1_IN_8 => UNWINDOWED_227 ,
										MUX_10_1_IN_9 => UNWINDOWED_738 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_369
									);
MUX_REORD_UNIT_370 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_370 ,
										MUX_10_1_IN_1 => UNWINDOWED_369 ,
										MUX_10_1_IN_2 => UNWINDOWED_372 ,
										MUX_10_1_IN_3 => UNWINDOWED_372 ,
										MUX_10_1_IN_4 => UNWINDOWED_357 ,
										MUX_10_1_IN_5 => UNWINDOWED_357 ,
										MUX_10_1_IN_6 => UNWINDOWED_357 ,
										MUX_10_1_IN_7 => UNWINDOWED_484 ,
										MUX_10_1_IN_8 => UNWINDOWED_229 ,
										MUX_10_1_IN_9 => UNWINDOWED_740 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_370
									);
MUX_REORD_UNIT_371 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_371 ,
										MUX_10_1_IN_1 => UNWINDOWED_371 ,
										MUX_10_1_IN_2 => UNWINDOWED_374 ,
										MUX_10_1_IN_3 => UNWINDOWED_374 ,
										MUX_10_1_IN_4 => UNWINDOWED_359 ,
										MUX_10_1_IN_5 => UNWINDOWED_359 ,
										MUX_10_1_IN_6 => UNWINDOWED_359 ,
										MUX_10_1_IN_7 => UNWINDOWED_486 ,
										MUX_10_1_IN_8 => UNWINDOWED_231 ,
										MUX_10_1_IN_9 => UNWINDOWED_742 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_371
									);
MUX_REORD_UNIT_372 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_372 ,
										MUX_10_1_IN_1 => UNWINDOWED_372 ,
										MUX_10_1_IN_2 => UNWINDOWED_369 ,
										MUX_10_1_IN_3 => UNWINDOWED_376 ,
										MUX_10_1_IN_4 => UNWINDOWED_361 ,
										MUX_10_1_IN_5 => UNWINDOWED_361 ,
										MUX_10_1_IN_6 => UNWINDOWED_361 ,
										MUX_10_1_IN_7 => UNWINDOWED_488 ,
										MUX_10_1_IN_8 => UNWINDOWED_233 ,
										MUX_10_1_IN_9 => UNWINDOWED_744 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_372
									);
MUX_REORD_UNIT_373 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_373 ,
										MUX_10_1_IN_1 => UNWINDOWED_374 ,
										MUX_10_1_IN_2 => UNWINDOWED_371 ,
										MUX_10_1_IN_3 => UNWINDOWED_378 ,
										MUX_10_1_IN_4 => UNWINDOWED_363 ,
										MUX_10_1_IN_5 => UNWINDOWED_363 ,
										MUX_10_1_IN_6 => UNWINDOWED_363 ,
										MUX_10_1_IN_7 => UNWINDOWED_490 ,
										MUX_10_1_IN_8 => UNWINDOWED_235 ,
										MUX_10_1_IN_9 => UNWINDOWED_746 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_373
									);
MUX_REORD_UNIT_374 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_374 ,
										MUX_10_1_IN_1 => UNWINDOWED_373 ,
										MUX_10_1_IN_2 => UNWINDOWED_373 ,
										MUX_10_1_IN_3 => UNWINDOWED_380 ,
										MUX_10_1_IN_4 => UNWINDOWED_365 ,
										MUX_10_1_IN_5 => UNWINDOWED_365 ,
										MUX_10_1_IN_6 => UNWINDOWED_365 ,
										MUX_10_1_IN_7 => UNWINDOWED_492 ,
										MUX_10_1_IN_8 => UNWINDOWED_237 ,
										MUX_10_1_IN_9 => UNWINDOWED_748 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_374
									);
MUX_REORD_UNIT_375 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_375 ,
										MUX_10_1_IN_1 => UNWINDOWED_375 ,
										MUX_10_1_IN_2 => UNWINDOWED_375 ,
										MUX_10_1_IN_3 => UNWINDOWED_382 ,
										MUX_10_1_IN_4 => UNWINDOWED_367 ,
										MUX_10_1_IN_5 => UNWINDOWED_367 ,
										MUX_10_1_IN_6 => UNWINDOWED_367 ,
										MUX_10_1_IN_7 => UNWINDOWED_494 ,
										MUX_10_1_IN_8 => UNWINDOWED_239 ,
										MUX_10_1_IN_9 => UNWINDOWED_750 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_375
									);
MUX_REORD_UNIT_376 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_376 ,
										MUX_10_1_IN_1 => UNWINDOWED_376 ,
										MUX_10_1_IN_2 => UNWINDOWED_376 ,
										MUX_10_1_IN_3 => UNWINDOWED_369 ,
										MUX_10_1_IN_4 => UNWINDOWED_369 ,
										MUX_10_1_IN_5 => UNWINDOWED_369 ,
										MUX_10_1_IN_6 => UNWINDOWED_369 ,
										MUX_10_1_IN_7 => UNWINDOWED_496 ,
										MUX_10_1_IN_8 => UNWINDOWED_241 ,
										MUX_10_1_IN_9 => UNWINDOWED_752 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_376
									);
MUX_REORD_UNIT_377 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_377 ,
										MUX_10_1_IN_1 => UNWINDOWED_378 ,
										MUX_10_1_IN_2 => UNWINDOWED_378 ,
										MUX_10_1_IN_3 => UNWINDOWED_371 ,
										MUX_10_1_IN_4 => UNWINDOWED_371 ,
										MUX_10_1_IN_5 => UNWINDOWED_371 ,
										MUX_10_1_IN_6 => UNWINDOWED_371 ,
										MUX_10_1_IN_7 => UNWINDOWED_498 ,
										MUX_10_1_IN_8 => UNWINDOWED_243 ,
										MUX_10_1_IN_9 => UNWINDOWED_754 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_377
									);
MUX_REORD_UNIT_378 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_378 ,
										MUX_10_1_IN_1 => UNWINDOWED_377 ,
										MUX_10_1_IN_2 => UNWINDOWED_380 ,
										MUX_10_1_IN_3 => UNWINDOWED_373 ,
										MUX_10_1_IN_4 => UNWINDOWED_373 ,
										MUX_10_1_IN_5 => UNWINDOWED_373 ,
										MUX_10_1_IN_6 => UNWINDOWED_373 ,
										MUX_10_1_IN_7 => UNWINDOWED_500 ,
										MUX_10_1_IN_8 => UNWINDOWED_245 ,
										MUX_10_1_IN_9 => UNWINDOWED_756 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_378
									);
MUX_REORD_UNIT_379 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_379 ,
										MUX_10_1_IN_1 => UNWINDOWED_379 ,
										MUX_10_1_IN_2 => UNWINDOWED_382 ,
										MUX_10_1_IN_3 => UNWINDOWED_375 ,
										MUX_10_1_IN_4 => UNWINDOWED_375 ,
										MUX_10_1_IN_5 => UNWINDOWED_375 ,
										MUX_10_1_IN_6 => UNWINDOWED_375 ,
										MUX_10_1_IN_7 => UNWINDOWED_502 ,
										MUX_10_1_IN_8 => UNWINDOWED_247 ,
										MUX_10_1_IN_9 => UNWINDOWED_758 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_379
									);
MUX_REORD_UNIT_380 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_380 ,
										MUX_10_1_IN_1 => UNWINDOWED_380 ,
										MUX_10_1_IN_2 => UNWINDOWED_377 ,
										MUX_10_1_IN_3 => UNWINDOWED_377 ,
										MUX_10_1_IN_4 => UNWINDOWED_377 ,
										MUX_10_1_IN_5 => UNWINDOWED_377 ,
										MUX_10_1_IN_6 => UNWINDOWED_377 ,
										MUX_10_1_IN_7 => UNWINDOWED_504 ,
										MUX_10_1_IN_8 => UNWINDOWED_249 ,
										MUX_10_1_IN_9 => UNWINDOWED_760 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_380
									);
MUX_REORD_UNIT_381 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_381 ,
										MUX_10_1_IN_1 => UNWINDOWED_382 ,
										MUX_10_1_IN_2 => UNWINDOWED_379 ,
										MUX_10_1_IN_3 => UNWINDOWED_379 ,
										MUX_10_1_IN_4 => UNWINDOWED_379 ,
										MUX_10_1_IN_5 => UNWINDOWED_379 ,
										MUX_10_1_IN_6 => UNWINDOWED_379 ,
										MUX_10_1_IN_7 => UNWINDOWED_506 ,
										MUX_10_1_IN_8 => UNWINDOWED_251 ,
										MUX_10_1_IN_9 => UNWINDOWED_762 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_381
									);
MUX_REORD_UNIT_382 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_382 ,
										MUX_10_1_IN_1 => UNWINDOWED_381 ,
										MUX_10_1_IN_2 => UNWINDOWED_381 ,
										MUX_10_1_IN_3 => UNWINDOWED_381 ,
										MUX_10_1_IN_4 => UNWINDOWED_381 ,
										MUX_10_1_IN_5 => UNWINDOWED_381 ,
										MUX_10_1_IN_6 => UNWINDOWED_381 ,
										MUX_10_1_IN_7 => UNWINDOWED_508 ,
										MUX_10_1_IN_8 => UNWINDOWED_253 ,
										MUX_10_1_IN_9 => UNWINDOWED_764 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_382
									);
MUX_REORD_UNIT_383 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_383 ,
										MUX_10_1_IN_1 => UNWINDOWED_383 ,
										MUX_10_1_IN_2 => UNWINDOWED_383 ,
										MUX_10_1_IN_3 => UNWINDOWED_383 ,
										MUX_10_1_IN_4 => UNWINDOWED_383 ,
										MUX_10_1_IN_5 => UNWINDOWED_383 ,
										MUX_10_1_IN_6 => UNWINDOWED_383 ,
										MUX_10_1_IN_7 => UNWINDOWED_510 ,
										MUX_10_1_IN_8 => UNWINDOWED_255 ,
										MUX_10_1_IN_9 => UNWINDOWED_766 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_383
									);
MUX_REORD_UNIT_384 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_384 ,
										MUX_10_1_IN_1 => UNWINDOWED_384 ,
										MUX_10_1_IN_2 => UNWINDOWED_384 ,
										MUX_10_1_IN_3 => UNWINDOWED_384 ,
										MUX_10_1_IN_4 => UNWINDOWED_384 ,
										MUX_10_1_IN_5 => UNWINDOWED_384 ,
										MUX_10_1_IN_6 => UNWINDOWED_384 ,
										MUX_10_1_IN_7 => UNWINDOWED_257 ,
										MUX_10_1_IN_8 => UNWINDOWED_257 ,
										MUX_10_1_IN_9 => UNWINDOWED_768 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_384
									);
MUX_REORD_UNIT_385 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_385 ,
										MUX_10_1_IN_1 => UNWINDOWED_386 ,
										MUX_10_1_IN_2 => UNWINDOWED_386 ,
										MUX_10_1_IN_3 => UNWINDOWED_386 ,
										MUX_10_1_IN_4 => UNWINDOWED_386 ,
										MUX_10_1_IN_5 => UNWINDOWED_386 ,
										MUX_10_1_IN_6 => UNWINDOWED_386 ,
										MUX_10_1_IN_7 => UNWINDOWED_259 ,
										MUX_10_1_IN_8 => UNWINDOWED_259 ,
										MUX_10_1_IN_9 => UNWINDOWED_770 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_385
									);
MUX_REORD_UNIT_386 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_386 ,
										MUX_10_1_IN_1 => UNWINDOWED_385 ,
										MUX_10_1_IN_2 => UNWINDOWED_388 ,
										MUX_10_1_IN_3 => UNWINDOWED_388 ,
										MUX_10_1_IN_4 => UNWINDOWED_388 ,
										MUX_10_1_IN_5 => UNWINDOWED_388 ,
										MUX_10_1_IN_6 => UNWINDOWED_388 ,
										MUX_10_1_IN_7 => UNWINDOWED_261 ,
										MUX_10_1_IN_8 => UNWINDOWED_261 ,
										MUX_10_1_IN_9 => UNWINDOWED_772 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_386
									);
MUX_REORD_UNIT_387 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_387 ,
										MUX_10_1_IN_1 => UNWINDOWED_387 ,
										MUX_10_1_IN_2 => UNWINDOWED_390 ,
										MUX_10_1_IN_3 => UNWINDOWED_390 ,
										MUX_10_1_IN_4 => UNWINDOWED_390 ,
										MUX_10_1_IN_5 => UNWINDOWED_390 ,
										MUX_10_1_IN_6 => UNWINDOWED_390 ,
										MUX_10_1_IN_7 => UNWINDOWED_263 ,
										MUX_10_1_IN_8 => UNWINDOWED_263 ,
										MUX_10_1_IN_9 => UNWINDOWED_774 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_387
									);
MUX_REORD_UNIT_388 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_388 ,
										MUX_10_1_IN_1 => UNWINDOWED_388 ,
										MUX_10_1_IN_2 => UNWINDOWED_385 ,
										MUX_10_1_IN_3 => UNWINDOWED_392 ,
										MUX_10_1_IN_4 => UNWINDOWED_392 ,
										MUX_10_1_IN_5 => UNWINDOWED_392 ,
										MUX_10_1_IN_6 => UNWINDOWED_392 ,
										MUX_10_1_IN_7 => UNWINDOWED_265 ,
										MUX_10_1_IN_8 => UNWINDOWED_265 ,
										MUX_10_1_IN_9 => UNWINDOWED_776 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_388
									);
MUX_REORD_UNIT_389 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_389 ,
										MUX_10_1_IN_1 => UNWINDOWED_390 ,
										MUX_10_1_IN_2 => UNWINDOWED_387 ,
										MUX_10_1_IN_3 => UNWINDOWED_394 ,
										MUX_10_1_IN_4 => UNWINDOWED_394 ,
										MUX_10_1_IN_5 => UNWINDOWED_394 ,
										MUX_10_1_IN_6 => UNWINDOWED_394 ,
										MUX_10_1_IN_7 => UNWINDOWED_267 ,
										MUX_10_1_IN_8 => UNWINDOWED_267 ,
										MUX_10_1_IN_9 => UNWINDOWED_778 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_389
									);
MUX_REORD_UNIT_390 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_390 ,
										MUX_10_1_IN_1 => UNWINDOWED_389 ,
										MUX_10_1_IN_2 => UNWINDOWED_389 ,
										MUX_10_1_IN_3 => UNWINDOWED_396 ,
										MUX_10_1_IN_4 => UNWINDOWED_396 ,
										MUX_10_1_IN_5 => UNWINDOWED_396 ,
										MUX_10_1_IN_6 => UNWINDOWED_396 ,
										MUX_10_1_IN_7 => UNWINDOWED_269 ,
										MUX_10_1_IN_8 => UNWINDOWED_269 ,
										MUX_10_1_IN_9 => UNWINDOWED_780 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_390
									);
MUX_REORD_UNIT_391 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_391 ,
										MUX_10_1_IN_1 => UNWINDOWED_391 ,
										MUX_10_1_IN_2 => UNWINDOWED_391 ,
										MUX_10_1_IN_3 => UNWINDOWED_398 ,
										MUX_10_1_IN_4 => UNWINDOWED_398 ,
										MUX_10_1_IN_5 => UNWINDOWED_398 ,
										MUX_10_1_IN_6 => UNWINDOWED_398 ,
										MUX_10_1_IN_7 => UNWINDOWED_271 ,
										MUX_10_1_IN_8 => UNWINDOWED_271 ,
										MUX_10_1_IN_9 => UNWINDOWED_782 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_391
									);
MUX_REORD_UNIT_392 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_392 ,
										MUX_10_1_IN_1 => UNWINDOWED_392 ,
										MUX_10_1_IN_2 => UNWINDOWED_392 ,
										MUX_10_1_IN_3 => UNWINDOWED_385 ,
										MUX_10_1_IN_4 => UNWINDOWED_400 ,
										MUX_10_1_IN_5 => UNWINDOWED_400 ,
										MUX_10_1_IN_6 => UNWINDOWED_400 ,
										MUX_10_1_IN_7 => UNWINDOWED_273 ,
										MUX_10_1_IN_8 => UNWINDOWED_273 ,
										MUX_10_1_IN_9 => UNWINDOWED_784 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_392
									);
MUX_REORD_UNIT_393 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_393 ,
										MUX_10_1_IN_1 => UNWINDOWED_394 ,
										MUX_10_1_IN_2 => UNWINDOWED_394 ,
										MUX_10_1_IN_3 => UNWINDOWED_387 ,
										MUX_10_1_IN_4 => UNWINDOWED_402 ,
										MUX_10_1_IN_5 => UNWINDOWED_402 ,
										MUX_10_1_IN_6 => UNWINDOWED_402 ,
										MUX_10_1_IN_7 => UNWINDOWED_275 ,
										MUX_10_1_IN_8 => UNWINDOWED_275 ,
										MUX_10_1_IN_9 => UNWINDOWED_786 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_393
									);
MUX_REORD_UNIT_394 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_394 ,
										MUX_10_1_IN_1 => UNWINDOWED_393 ,
										MUX_10_1_IN_2 => UNWINDOWED_396 ,
										MUX_10_1_IN_3 => UNWINDOWED_389 ,
										MUX_10_1_IN_4 => UNWINDOWED_404 ,
										MUX_10_1_IN_5 => UNWINDOWED_404 ,
										MUX_10_1_IN_6 => UNWINDOWED_404 ,
										MUX_10_1_IN_7 => UNWINDOWED_277 ,
										MUX_10_1_IN_8 => UNWINDOWED_277 ,
										MUX_10_1_IN_9 => UNWINDOWED_788 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_394
									);
MUX_REORD_UNIT_395 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_395 ,
										MUX_10_1_IN_1 => UNWINDOWED_395 ,
										MUX_10_1_IN_2 => UNWINDOWED_398 ,
										MUX_10_1_IN_3 => UNWINDOWED_391 ,
										MUX_10_1_IN_4 => UNWINDOWED_406 ,
										MUX_10_1_IN_5 => UNWINDOWED_406 ,
										MUX_10_1_IN_6 => UNWINDOWED_406 ,
										MUX_10_1_IN_7 => UNWINDOWED_279 ,
										MUX_10_1_IN_8 => UNWINDOWED_279 ,
										MUX_10_1_IN_9 => UNWINDOWED_790 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_395
									);
MUX_REORD_UNIT_396 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_396 ,
										MUX_10_1_IN_1 => UNWINDOWED_396 ,
										MUX_10_1_IN_2 => UNWINDOWED_393 ,
										MUX_10_1_IN_3 => UNWINDOWED_393 ,
										MUX_10_1_IN_4 => UNWINDOWED_408 ,
										MUX_10_1_IN_5 => UNWINDOWED_408 ,
										MUX_10_1_IN_6 => UNWINDOWED_408 ,
										MUX_10_1_IN_7 => UNWINDOWED_281 ,
										MUX_10_1_IN_8 => UNWINDOWED_281 ,
										MUX_10_1_IN_9 => UNWINDOWED_792 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_396
									);
MUX_REORD_UNIT_397 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_397 ,
										MUX_10_1_IN_1 => UNWINDOWED_398 ,
										MUX_10_1_IN_2 => UNWINDOWED_395 ,
										MUX_10_1_IN_3 => UNWINDOWED_395 ,
										MUX_10_1_IN_4 => UNWINDOWED_410 ,
										MUX_10_1_IN_5 => UNWINDOWED_410 ,
										MUX_10_1_IN_6 => UNWINDOWED_410 ,
										MUX_10_1_IN_7 => UNWINDOWED_283 ,
										MUX_10_1_IN_8 => UNWINDOWED_283 ,
										MUX_10_1_IN_9 => UNWINDOWED_794 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_397
									);
MUX_REORD_UNIT_398 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_398 ,
										MUX_10_1_IN_1 => UNWINDOWED_397 ,
										MUX_10_1_IN_2 => UNWINDOWED_397 ,
										MUX_10_1_IN_3 => UNWINDOWED_397 ,
										MUX_10_1_IN_4 => UNWINDOWED_412 ,
										MUX_10_1_IN_5 => UNWINDOWED_412 ,
										MUX_10_1_IN_6 => UNWINDOWED_412 ,
										MUX_10_1_IN_7 => UNWINDOWED_285 ,
										MUX_10_1_IN_8 => UNWINDOWED_285 ,
										MUX_10_1_IN_9 => UNWINDOWED_796 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_398
									);
MUX_REORD_UNIT_399 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_399 ,
										MUX_10_1_IN_1 => UNWINDOWED_399 ,
										MUX_10_1_IN_2 => UNWINDOWED_399 ,
										MUX_10_1_IN_3 => UNWINDOWED_399 ,
										MUX_10_1_IN_4 => UNWINDOWED_414 ,
										MUX_10_1_IN_5 => UNWINDOWED_414 ,
										MUX_10_1_IN_6 => UNWINDOWED_414 ,
										MUX_10_1_IN_7 => UNWINDOWED_287 ,
										MUX_10_1_IN_8 => UNWINDOWED_287 ,
										MUX_10_1_IN_9 => UNWINDOWED_798 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_399
									);
MUX_REORD_UNIT_400 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_400 ,
										MUX_10_1_IN_1 => UNWINDOWED_400 ,
										MUX_10_1_IN_2 => UNWINDOWED_400 ,
										MUX_10_1_IN_3 => UNWINDOWED_400 ,
										MUX_10_1_IN_4 => UNWINDOWED_385 ,
										MUX_10_1_IN_5 => UNWINDOWED_416 ,
										MUX_10_1_IN_6 => UNWINDOWED_416 ,
										MUX_10_1_IN_7 => UNWINDOWED_289 ,
										MUX_10_1_IN_8 => UNWINDOWED_289 ,
										MUX_10_1_IN_9 => UNWINDOWED_800 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_400
									);
MUX_REORD_UNIT_401 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_401 ,
										MUX_10_1_IN_1 => UNWINDOWED_402 ,
										MUX_10_1_IN_2 => UNWINDOWED_402 ,
										MUX_10_1_IN_3 => UNWINDOWED_402 ,
										MUX_10_1_IN_4 => UNWINDOWED_387 ,
										MUX_10_1_IN_5 => UNWINDOWED_418 ,
										MUX_10_1_IN_6 => UNWINDOWED_418 ,
										MUX_10_1_IN_7 => UNWINDOWED_291 ,
										MUX_10_1_IN_8 => UNWINDOWED_291 ,
										MUX_10_1_IN_9 => UNWINDOWED_802 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_401
									);
MUX_REORD_UNIT_402 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_402 ,
										MUX_10_1_IN_1 => UNWINDOWED_401 ,
										MUX_10_1_IN_2 => UNWINDOWED_404 ,
										MUX_10_1_IN_3 => UNWINDOWED_404 ,
										MUX_10_1_IN_4 => UNWINDOWED_389 ,
										MUX_10_1_IN_5 => UNWINDOWED_420 ,
										MUX_10_1_IN_6 => UNWINDOWED_420 ,
										MUX_10_1_IN_7 => UNWINDOWED_293 ,
										MUX_10_1_IN_8 => UNWINDOWED_293 ,
										MUX_10_1_IN_9 => UNWINDOWED_804 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_402
									);
MUX_REORD_UNIT_403 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_403 ,
										MUX_10_1_IN_1 => UNWINDOWED_403 ,
										MUX_10_1_IN_2 => UNWINDOWED_406 ,
										MUX_10_1_IN_3 => UNWINDOWED_406 ,
										MUX_10_1_IN_4 => UNWINDOWED_391 ,
										MUX_10_1_IN_5 => UNWINDOWED_422 ,
										MUX_10_1_IN_6 => UNWINDOWED_422 ,
										MUX_10_1_IN_7 => UNWINDOWED_295 ,
										MUX_10_1_IN_8 => UNWINDOWED_295 ,
										MUX_10_1_IN_9 => UNWINDOWED_806 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_403
									);
MUX_REORD_UNIT_404 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_404 ,
										MUX_10_1_IN_1 => UNWINDOWED_404 ,
										MUX_10_1_IN_2 => UNWINDOWED_401 ,
										MUX_10_1_IN_3 => UNWINDOWED_408 ,
										MUX_10_1_IN_4 => UNWINDOWED_393 ,
										MUX_10_1_IN_5 => UNWINDOWED_424 ,
										MUX_10_1_IN_6 => UNWINDOWED_424 ,
										MUX_10_1_IN_7 => UNWINDOWED_297 ,
										MUX_10_1_IN_8 => UNWINDOWED_297 ,
										MUX_10_1_IN_9 => UNWINDOWED_808 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_404
									);
MUX_REORD_UNIT_405 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_405 ,
										MUX_10_1_IN_1 => UNWINDOWED_406 ,
										MUX_10_1_IN_2 => UNWINDOWED_403 ,
										MUX_10_1_IN_3 => UNWINDOWED_410 ,
										MUX_10_1_IN_4 => UNWINDOWED_395 ,
										MUX_10_1_IN_5 => UNWINDOWED_426 ,
										MUX_10_1_IN_6 => UNWINDOWED_426 ,
										MUX_10_1_IN_7 => UNWINDOWED_299 ,
										MUX_10_1_IN_8 => UNWINDOWED_299 ,
										MUX_10_1_IN_9 => UNWINDOWED_810 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_405
									);
MUX_REORD_UNIT_406 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_406 ,
										MUX_10_1_IN_1 => UNWINDOWED_405 ,
										MUX_10_1_IN_2 => UNWINDOWED_405 ,
										MUX_10_1_IN_3 => UNWINDOWED_412 ,
										MUX_10_1_IN_4 => UNWINDOWED_397 ,
										MUX_10_1_IN_5 => UNWINDOWED_428 ,
										MUX_10_1_IN_6 => UNWINDOWED_428 ,
										MUX_10_1_IN_7 => UNWINDOWED_301 ,
										MUX_10_1_IN_8 => UNWINDOWED_301 ,
										MUX_10_1_IN_9 => UNWINDOWED_812 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_406
									);
MUX_REORD_UNIT_407 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_407 ,
										MUX_10_1_IN_1 => UNWINDOWED_407 ,
										MUX_10_1_IN_2 => UNWINDOWED_407 ,
										MUX_10_1_IN_3 => UNWINDOWED_414 ,
										MUX_10_1_IN_4 => UNWINDOWED_399 ,
										MUX_10_1_IN_5 => UNWINDOWED_430 ,
										MUX_10_1_IN_6 => UNWINDOWED_430 ,
										MUX_10_1_IN_7 => UNWINDOWED_303 ,
										MUX_10_1_IN_8 => UNWINDOWED_303 ,
										MUX_10_1_IN_9 => UNWINDOWED_814 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_407
									);
MUX_REORD_UNIT_408 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_408 ,
										MUX_10_1_IN_1 => UNWINDOWED_408 ,
										MUX_10_1_IN_2 => UNWINDOWED_408 ,
										MUX_10_1_IN_3 => UNWINDOWED_401 ,
										MUX_10_1_IN_4 => UNWINDOWED_401 ,
										MUX_10_1_IN_5 => UNWINDOWED_432 ,
										MUX_10_1_IN_6 => UNWINDOWED_432 ,
										MUX_10_1_IN_7 => UNWINDOWED_305 ,
										MUX_10_1_IN_8 => UNWINDOWED_305 ,
										MUX_10_1_IN_9 => UNWINDOWED_816 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_408
									);
MUX_REORD_UNIT_409 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_409 ,
										MUX_10_1_IN_1 => UNWINDOWED_410 ,
										MUX_10_1_IN_2 => UNWINDOWED_410 ,
										MUX_10_1_IN_3 => UNWINDOWED_403 ,
										MUX_10_1_IN_4 => UNWINDOWED_403 ,
										MUX_10_1_IN_5 => UNWINDOWED_434 ,
										MUX_10_1_IN_6 => UNWINDOWED_434 ,
										MUX_10_1_IN_7 => UNWINDOWED_307 ,
										MUX_10_1_IN_8 => UNWINDOWED_307 ,
										MUX_10_1_IN_9 => UNWINDOWED_818 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_409
									);
MUX_REORD_UNIT_410 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_410 ,
										MUX_10_1_IN_1 => UNWINDOWED_409 ,
										MUX_10_1_IN_2 => UNWINDOWED_412 ,
										MUX_10_1_IN_3 => UNWINDOWED_405 ,
										MUX_10_1_IN_4 => UNWINDOWED_405 ,
										MUX_10_1_IN_5 => UNWINDOWED_436 ,
										MUX_10_1_IN_6 => UNWINDOWED_436 ,
										MUX_10_1_IN_7 => UNWINDOWED_309 ,
										MUX_10_1_IN_8 => UNWINDOWED_309 ,
										MUX_10_1_IN_9 => UNWINDOWED_820 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_410
									);
MUX_REORD_UNIT_411 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_411 ,
										MUX_10_1_IN_1 => UNWINDOWED_411 ,
										MUX_10_1_IN_2 => UNWINDOWED_414 ,
										MUX_10_1_IN_3 => UNWINDOWED_407 ,
										MUX_10_1_IN_4 => UNWINDOWED_407 ,
										MUX_10_1_IN_5 => UNWINDOWED_438 ,
										MUX_10_1_IN_6 => UNWINDOWED_438 ,
										MUX_10_1_IN_7 => UNWINDOWED_311 ,
										MUX_10_1_IN_8 => UNWINDOWED_311 ,
										MUX_10_1_IN_9 => UNWINDOWED_822 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_411
									);
MUX_REORD_UNIT_412 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_412 ,
										MUX_10_1_IN_1 => UNWINDOWED_412 ,
										MUX_10_1_IN_2 => UNWINDOWED_409 ,
										MUX_10_1_IN_3 => UNWINDOWED_409 ,
										MUX_10_1_IN_4 => UNWINDOWED_409 ,
										MUX_10_1_IN_5 => UNWINDOWED_440 ,
										MUX_10_1_IN_6 => UNWINDOWED_440 ,
										MUX_10_1_IN_7 => UNWINDOWED_313 ,
										MUX_10_1_IN_8 => UNWINDOWED_313 ,
										MUX_10_1_IN_9 => UNWINDOWED_824 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_412
									);
MUX_REORD_UNIT_413 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_413 ,
										MUX_10_1_IN_1 => UNWINDOWED_414 ,
										MUX_10_1_IN_2 => UNWINDOWED_411 ,
										MUX_10_1_IN_3 => UNWINDOWED_411 ,
										MUX_10_1_IN_4 => UNWINDOWED_411 ,
										MUX_10_1_IN_5 => UNWINDOWED_442 ,
										MUX_10_1_IN_6 => UNWINDOWED_442 ,
										MUX_10_1_IN_7 => UNWINDOWED_315 ,
										MUX_10_1_IN_8 => UNWINDOWED_315 ,
										MUX_10_1_IN_9 => UNWINDOWED_826 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_413
									);
MUX_REORD_UNIT_414 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_414 ,
										MUX_10_1_IN_1 => UNWINDOWED_413 ,
										MUX_10_1_IN_2 => UNWINDOWED_413 ,
										MUX_10_1_IN_3 => UNWINDOWED_413 ,
										MUX_10_1_IN_4 => UNWINDOWED_413 ,
										MUX_10_1_IN_5 => UNWINDOWED_444 ,
										MUX_10_1_IN_6 => UNWINDOWED_444 ,
										MUX_10_1_IN_7 => UNWINDOWED_317 ,
										MUX_10_1_IN_8 => UNWINDOWED_317 ,
										MUX_10_1_IN_9 => UNWINDOWED_828 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_414
									);
MUX_REORD_UNIT_415 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_415 ,
										MUX_10_1_IN_1 => UNWINDOWED_415 ,
										MUX_10_1_IN_2 => UNWINDOWED_415 ,
										MUX_10_1_IN_3 => UNWINDOWED_415 ,
										MUX_10_1_IN_4 => UNWINDOWED_415 ,
										MUX_10_1_IN_5 => UNWINDOWED_446 ,
										MUX_10_1_IN_6 => UNWINDOWED_446 ,
										MUX_10_1_IN_7 => UNWINDOWED_319 ,
										MUX_10_1_IN_8 => UNWINDOWED_319 ,
										MUX_10_1_IN_9 => UNWINDOWED_830 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_415
									);
MUX_REORD_UNIT_416 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_416 ,
										MUX_10_1_IN_1 => UNWINDOWED_416 ,
										MUX_10_1_IN_2 => UNWINDOWED_416 ,
										MUX_10_1_IN_3 => UNWINDOWED_416 ,
										MUX_10_1_IN_4 => UNWINDOWED_416 ,
										MUX_10_1_IN_5 => UNWINDOWED_385 ,
										MUX_10_1_IN_6 => UNWINDOWED_448 ,
										MUX_10_1_IN_7 => UNWINDOWED_321 ,
										MUX_10_1_IN_8 => UNWINDOWED_321 ,
										MUX_10_1_IN_9 => UNWINDOWED_832 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_416
									);
MUX_REORD_UNIT_417 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_417 ,
										MUX_10_1_IN_1 => UNWINDOWED_418 ,
										MUX_10_1_IN_2 => UNWINDOWED_418 ,
										MUX_10_1_IN_3 => UNWINDOWED_418 ,
										MUX_10_1_IN_4 => UNWINDOWED_418 ,
										MUX_10_1_IN_5 => UNWINDOWED_387 ,
										MUX_10_1_IN_6 => UNWINDOWED_450 ,
										MUX_10_1_IN_7 => UNWINDOWED_323 ,
										MUX_10_1_IN_8 => UNWINDOWED_323 ,
										MUX_10_1_IN_9 => UNWINDOWED_834 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_417
									);
MUX_REORD_UNIT_418 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_418 ,
										MUX_10_1_IN_1 => UNWINDOWED_417 ,
										MUX_10_1_IN_2 => UNWINDOWED_420 ,
										MUX_10_1_IN_3 => UNWINDOWED_420 ,
										MUX_10_1_IN_4 => UNWINDOWED_420 ,
										MUX_10_1_IN_5 => UNWINDOWED_389 ,
										MUX_10_1_IN_6 => UNWINDOWED_452 ,
										MUX_10_1_IN_7 => UNWINDOWED_325 ,
										MUX_10_1_IN_8 => UNWINDOWED_325 ,
										MUX_10_1_IN_9 => UNWINDOWED_836 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_418
									);
MUX_REORD_UNIT_419 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_419 ,
										MUX_10_1_IN_1 => UNWINDOWED_419 ,
										MUX_10_1_IN_2 => UNWINDOWED_422 ,
										MUX_10_1_IN_3 => UNWINDOWED_422 ,
										MUX_10_1_IN_4 => UNWINDOWED_422 ,
										MUX_10_1_IN_5 => UNWINDOWED_391 ,
										MUX_10_1_IN_6 => UNWINDOWED_454 ,
										MUX_10_1_IN_7 => UNWINDOWED_327 ,
										MUX_10_1_IN_8 => UNWINDOWED_327 ,
										MUX_10_1_IN_9 => UNWINDOWED_838 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_419
									);
MUX_REORD_UNIT_420 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_420 ,
										MUX_10_1_IN_1 => UNWINDOWED_420 ,
										MUX_10_1_IN_2 => UNWINDOWED_417 ,
										MUX_10_1_IN_3 => UNWINDOWED_424 ,
										MUX_10_1_IN_4 => UNWINDOWED_424 ,
										MUX_10_1_IN_5 => UNWINDOWED_393 ,
										MUX_10_1_IN_6 => UNWINDOWED_456 ,
										MUX_10_1_IN_7 => UNWINDOWED_329 ,
										MUX_10_1_IN_8 => UNWINDOWED_329 ,
										MUX_10_1_IN_9 => UNWINDOWED_840 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_420
									);
MUX_REORD_UNIT_421 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_421 ,
										MUX_10_1_IN_1 => UNWINDOWED_422 ,
										MUX_10_1_IN_2 => UNWINDOWED_419 ,
										MUX_10_1_IN_3 => UNWINDOWED_426 ,
										MUX_10_1_IN_4 => UNWINDOWED_426 ,
										MUX_10_1_IN_5 => UNWINDOWED_395 ,
										MUX_10_1_IN_6 => UNWINDOWED_458 ,
										MUX_10_1_IN_7 => UNWINDOWED_331 ,
										MUX_10_1_IN_8 => UNWINDOWED_331 ,
										MUX_10_1_IN_9 => UNWINDOWED_842 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_421
									);
MUX_REORD_UNIT_422 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_422 ,
										MUX_10_1_IN_1 => UNWINDOWED_421 ,
										MUX_10_1_IN_2 => UNWINDOWED_421 ,
										MUX_10_1_IN_3 => UNWINDOWED_428 ,
										MUX_10_1_IN_4 => UNWINDOWED_428 ,
										MUX_10_1_IN_5 => UNWINDOWED_397 ,
										MUX_10_1_IN_6 => UNWINDOWED_460 ,
										MUX_10_1_IN_7 => UNWINDOWED_333 ,
										MUX_10_1_IN_8 => UNWINDOWED_333 ,
										MUX_10_1_IN_9 => UNWINDOWED_844 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_422
									);
MUX_REORD_UNIT_423 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_423 ,
										MUX_10_1_IN_1 => UNWINDOWED_423 ,
										MUX_10_1_IN_2 => UNWINDOWED_423 ,
										MUX_10_1_IN_3 => UNWINDOWED_430 ,
										MUX_10_1_IN_4 => UNWINDOWED_430 ,
										MUX_10_1_IN_5 => UNWINDOWED_399 ,
										MUX_10_1_IN_6 => UNWINDOWED_462 ,
										MUX_10_1_IN_7 => UNWINDOWED_335 ,
										MUX_10_1_IN_8 => UNWINDOWED_335 ,
										MUX_10_1_IN_9 => UNWINDOWED_846 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_423
									);
MUX_REORD_UNIT_424 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_424 ,
										MUX_10_1_IN_1 => UNWINDOWED_424 ,
										MUX_10_1_IN_2 => UNWINDOWED_424 ,
										MUX_10_1_IN_3 => UNWINDOWED_417 ,
										MUX_10_1_IN_4 => UNWINDOWED_432 ,
										MUX_10_1_IN_5 => UNWINDOWED_401 ,
										MUX_10_1_IN_6 => UNWINDOWED_464 ,
										MUX_10_1_IN_7 => UNWINDOWED_337 ,
										MUX_10_1_IN_8 => UNWINDOWED_337 ,
										MUX_10_1_IN_9 => UNWINDOWED_848 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_424
									);
MUX_REORD_UNIT_425 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_425 ,
										MUX_10_1_IN_1 => UNWINDOWED_426 ,
										MUX_10_1_IN_2 => UNWINDOWED_426 ,
										MUX_10_1_IN_3 => UNWINDOWED_419 ,
										MUX_10_1_IN_4 => UNWINDOWED_434 ,
										MUX_10_1_IN_5 => UNWINDOWED_403 ,
										MUX_10_1_IN_6 => UNWINDOWED_466 ,
										MUX_10_1_IN_7 => UNWINDOWED_339 ,
										MUX_10_1_IN_8 => UNWINDOWED_339 ,
										MUX_10_1_IN_9 => UNWINDOWED_850 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_425
									);
MUX_REORD_UNIT_426 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_426 ,
										MUX_10_1_IN_1 => UNWINDOWED_425 ,
										MUX_10_1_IN_2 => UNWINDOWED_428 ,
										MUX_10_1_IN_3 => UNWINDOWED_421 ,
										MUX_10_1_IN_4 => UNWINDOWED_436 ,
										MUX_10_1_IN_5 => UNWINDOWED_405 ,
										MUX_10_1_IN_6 => UNWINDOWED_468 ,
										MUX_10_1_IN_7 => UNWINDOWED_341 ,
										MUX_10_1_IN_8 => UNWINDOWED_341 ,
										MUX_10_1_IN_9 => UNWINDOWED_852 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_426
									);
MUX_REORD_UNIT_427 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_427 ,
										MUX_10_1_IN_1 => UNWINDOWED_427 ,
										MUX_10_1_IN_2 => UNWINDOWED_430 ,
										MUX_10_1_IN_3 => UNWINDOWED_423 ,
										MUX_10_1_IN_4 => UNWINDOWED_438 ,
										MUX_10_1_IN_5 => UNWINDOWED_407 ,
										MUX_10_1_IN_6 => UNWINDOWED_470 ,
										MUX_10_1_IN_7 => UNWINDOWED_343 ,
										MUX_10_1_IN_8 => UNWINDOWED_343 ,
										MUX_10_1_IN_9 => UNWINDOWED_854 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_427
									);
MUX_REORD_UNIT_428 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_428 ,
										MUX_10_1_IN_1 => UNWINDOWED_428 ,
										MUX_10_1_IN_2 => UNWINDOWED_425 ,
										MUX_10_1_IN_3 => UNWINDOWED_425 ,
										MUX_10_1_IN_4 => UNWINDOWED_440 ,
										MUX_10_1_IN_5 => UNWINDOWED_409 ,
										MUX_10_1_IN_6 => UNWINDOWED_472 ,
										MUX_10_1_IN_7 => UNWINDOWED_345 ,
										MUX_10_1_IN_8 => UNWINDOWED_345 ,
										MUX_10_1_IN_9 => UNWINDOWED_856 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_428
									);
MUX_REORD_UNIT_429 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_429 ,
										MUX_10_1_IN_1 => UNWINDOWED_430 ,
										MUX_10_1_IN_2 => UNWINDOWED_427 ,
										MUX_10_1_IN_3 => UNWINDOWED_427 ,
										MUX_10_1_IN_4 => UNWINDOWED_442 ,
										MUX_10_1_IN_5 => UNWINDOWED_411 ,
										MUX_10_1_IN_6 => UNWINDOWED_474 ,
										MUX_10_1_IN_7 => UNWINDOWED_347 ,
										MUX_10_1_IN_8 => UNWINDOWED_347 ,
										MUX_10_1_IN_9 => UNWINDOWED_858 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_429
									);
MUX_REORD_UNIT_430 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_430 ,
										MUX_10_1_IN_1 => UNWINDOWED_429 ,
										MUX_10_1_IN_2 => UNWINDOWED_429 ,
										MUX_10_1_IN_3 => UNWINDOWED_429 ,
										MUX_10_1_IN_4 => UNWINDOWED_444 ,
										MUX_10_1_IN_5 => UNWINDOWED_413 ,
										MUX_10_1_IN_6 => UNWINDOWED_476 ,
										MUX_10_1_IN_7 => UNWINDOWED_349 ,
										MUX_10_1_IN_8 => UNWINDOWED_349 ,
										MUX_10_1_IN_9 => UNWINDOWED_860 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_430
									);
MUX_REORD_UNIT_431 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_431 ,
										MUX_10_1_IN_1 => UNWINDOWED_431 ,
										MUX_10_1_IN_2 => UNWINDOWED_431 ,
										MUX_10_1_IN_3 => UNWINDOWED_431 ,
										MUX_10_1_IN_4 => UNWINDOWED_446 ,
										MUX_10_1_IN_5 => UNWINDOWED_415 ,
										MUX_10_1_IN_6 => UNWINDOWED_478 ,
										MUX_10_1_IN_7 => UNWINDOWED_351 ,
										MUX_10_1_IN_8 => UNWINDOWED_351 ,
										MUX_10_1_IN_9 => UNWINDOWED_862 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_431
									);
MUX_REORD_UNIT_432 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_432 ,
										MUX_10_1_IN_1 => UNWINDOWED_432 ,
										MUX_10_1_IN_2 => UNWINDOWED_432 ,
										MUX_10_1_IN_3 => UNWINDOWED_432 ,
										MUX_10_1_IN_4 => UNWINDOWED_417 ,
										MUX_10_1_IN_5 => UNWINDOWED_417 ,
										MUX_10_1_IN_6 => UNWINDOWED_480 ,
										MUX_10_1_IN_7 => UNWINDOWED_353 ,
										MUX_10_1_IN_8 => UNWINDOWED_353 ,
										MUX_10_1_IN_9 => UNWINDOWED_864 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_432
									);
MUX_REORD_UNIT_433 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_433 ,
										MUX_10_1_IN_1 => UNWINDOWED_434 ,
										MUX_10_1_IN_2 => UNWINDOWED_434 ,
										MUX_10_1_IN_3 => UNWINDOWED_434 ,
										MUX_10_1_IN_4 => UNWINDOWED_419 ,
										MUX_10_1_IN_5 => UNWINDOWED_419 ,
										MUX_10_1_IN_6 => UNWINDOWED_482 ,
										MUX_10_1_IN_7 => UNWINDOWED_355 ,
										MUX_10_1_IN_8 => UNWINDOWED_355 ,
										MUX_10_1_IN_9 => UNWINDOWED_866 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_433
									);
MUX_REORD_UNIT_434 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_434 ,
										MUX_10_1_IN_1 => UNWINDOWED_433 ,
										MUX_10_1_IN_2 => UNWINDOWED_436 ,
										MUX_10_1_IN_3 => UNWINDOWED_436 ,
										MUX_10_1_IN_4 => UNWINDOWED_421 ,
										MUX_10_1_IN_5 => UNWINDOWED_421 ,
										MUX_10_1_IN_6 => UNWINDOWED_484 ,
										MUX_10_1_IN_7 => UNWINDOWED_357 ,
										MUX_10_1_IN_8 => UNWINDOWED_357 ,
										MUX_10_1_IN_9 => UNWINDOWED_868 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_434
									);
MUX_REORD_UNIT_435 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_435 ,
										MUX_10_1_IN_1 => UNWINDOWED_435 ,
										MUX_10_1_IN_2 => UNWINDOWED_438 ,
										MUX_10_1_IN_3 => UNWINDOWED_438 ,
										MUX_10_1_IN_4 => UNWINDOWED_423 ,
										MUX_10_1_IN_5 => UNWINDOWED_423 ,
										MUX_10_1_IN_6 => UNWINDOWED_486 ,
										MUX_10_1_IN_7 => UNWINDOWED_359 ,
										MUX_10_1_IN_8 => UNWINDOWED_359 ,
										MUX_10_1_IN_9 => UNWINDOWED_870 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_435
									);
MUX_REORD_UNIT_436 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_436 ,
										MUX_10_1_IN_1 => UNWINDOWED_436 ,
										MUX_10_1_IN_2 => UNWINDOWED_433 ,
										MUX_10_1_IN_3 => UNWINDOWED_440 ,
										MUX_10_1_IN_4 => UNWINDOWED_425 ,
										MUX_10_1_IN_5 => UNWINDOWED_425 ,
										MUX_10_1_IN_6 => UNWINDOWED_488 ,
										MUX_10_1_IN_7 => UNWINDOWED_361 ,
										MUX_10_1_IN_8 => UNWINDOWED_361 ,
										MUX_10_1_IN_9 => UNWINDOWED_872 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_436
									);
MUX_REORD_UNIT_437 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_437 ,
										MUX_10_1_IN_1 => UNWINDOWED_438 ,
										MUX_10_1_IN_2 => UNWINDOWED_435 ,
										MUX_10_1_IN_3 => UNWINDOWED_442 ,
										MUX_10_1_IN_4 => UNWINDOWED_427 ,
										MUX_10_1_IN_5 => UNWINDOWED_427 ,
										MUX_10_1_IN_6 => UNWINDOWED_490 ,
										MUX_10_1_IN_7 => UNWINDOWED_363 ,
										MUX_10_1_IN_8 => UNWINDOWED_363 ,
										MUX_10_1_IN_9 => UNWINDOWED_874 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_437
									);
MUX_REORD_UNIT_438 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_438 ,
										MUX_10_1_IN_1 => UNWINDOWED_437 ,
										MUX_10_1_IN_2 => UNWINDOWED_437 ,
										MUX_10_1_IN_3 => UNWINDOWED_444 ,
										MUX_10_1_IN_4 => UNWINDOWED_429 ,
										MUX_10_1_IN_5 => UNWINDOWED_429 ,
										MUX_10_1_IN_6 => UNWINDOWED_492 ,
										MUX_10_1_IN_7 => UNWINDOWED_365 ,
										MUX_10_1_IN_8 => UNWINDOWED_365 ,
										MUX_10_1_IN_9 => UNWINDOWED_876 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_438
									);
MUX_REORD_UNIT_439 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_439 ,
										MUX_10_1_IN_1 => UNWINDOWED_439 ,
										MUX_10_1_IN_2 => UNWINDOWED_439 ,
										MUX_10_1_IN_3 => UNWINDOWED_446 ,
										MUX_10_1_IN_4 => UNWINDOWED_431 ,
										MUX_10_1_IN_5 => UNWINDOWED_431 ,
										MUX_10_1_IN_6 => UNWINDOWED_494 ,
										MUX_10_1_IN_7 => UNWINDOWED_367 ,
										MUX_10_1_IN_8 => UNWINDOWED_367 ,
										MUX_10_1_IN_9 => UNWINDOWED_878 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_439
									);
MUX_REORD_UNIT_440 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_440 ,
										MUX_10_1_IN_1 => UNWINDOWED_440 ,
										MUX_10_1_IN_2 => UNWINDOWED_440 ,
										MUX_10_1_IN_3 => UNWINDOWED_433 ,
										MUX_10_1_IN_4 => UNWINDOWED_433 ,
										MUX_10_1_IN_5 => UNWINDOWED_433 ,
										MUX_10_1_IN_6 => UNWINDOWED_496 ,
										MUX_10_1_IN_7 => UNWINDOWED_369 ,
										MUX_10_1_IN_8 => UNWINDOWED_369 ,
										MUX_10_1_IN_9 => UNWINDOWED_880 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_440
									);
MUX_REORD_UNIT_441 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_441 ,
										MUX_10_1_IN_1 => UNWINDOWED_442 ,
										MUX_10_1_IN_2 => UNWINDOWED_442 ,
										MUX_10_1_IN_3 => UNWINDOWED_435 ,
										MUX_10_1_IN_4 => UNWINDOWED_435 ,
										MUX_10_1_IN_5 => UNWINDOWED_435 ,
										MUX_10_1_IN_6 => UNWINDOWED_498 ,
										MUX_10_1_IN_7 => UNWINDOWED_371 ,
										MUX_10_1_IN_8 => UNWINDOWED_371 ,
										MUX_10_1_IN_9 => UNWINDOWED_882 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_441
									);
MUX_REORD_UNIT_442 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_442 ,
										MUX_10_1_IN_1 => UNWINDOWED_441 ,
										MUX_10_1_IN_2 => UNWINDOWED_444 ,
										MUX_10_1_IN_3 => UNWINDOWED_437 ,
										MUX_10_1_IN_4 => UNWINDOWED_437 ,
										MUX_10_1_IN_5 => UNWINDOWED_437 ,
										MUX_10_1_IN_6 => UNWINDOWED_500 ,
										MUX_10_1_IN_7 => UNWINDOWED_373 ,
										MUX_10_1_IN_8 => UNWINDOWED_373 ,
										MUX_10_1_IN_9 => UNWINDOWED_884 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_442
									);
MUX_REORD_UNIT_443 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_443 ,
										MUX_10_1_IN_1 => UNWINDOWED_443 ,
										MUX_10_1_IN_2 => UNWINDOWED_446 ,
										MUX_10_1_IN_3 => UNWINDOWED_439 ,
										MUX_10_1_IN_4 => UNWINDOWED_439 ,
										MUX_10_1_IN_5 => UNWINDOWED_439 ,
										MUX_10_1_IN_6 => UNWINDOWED_502 ,
										MUX_10_1_IN_7 => UNWINDOWED_375 ,
										MUX_10_1_IN_8 => UNWINDOWED_375 ,
										MUX_10_1_IN_9 => UNWINDOWED_886 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_443
									);
MUX_REORD_UNIT_444 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_444 ,
										MUX_10_1_IN_1 => UNWINDOWED_444 ,
										MUX_10_1_IN_2 => UNWINDOWED_441 ,
										MUX_10_1_IN_3 => UNWINDOWED_441 ,
										MUX_10_1_IN_4 => UNWINDOWED_441 ,
										MUX_10_1_IN_5 => UNWINDOWED_441 ,
										MUX_10_1_IN_6 => UNWINDOWED_504 ,
										MUX_10_1_IN_7 => UNWINDOWED_377 ,
										MUX_10_1_IN_8 => UNWINDOWED_377 ,
										MUX_10_1_IN_9 => UNWINDOWED_888 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_444
									);
MUX_REORD_UNIT_445 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_445 ,
										MUX_10_1_IN_1 => UNWINDOWED_446 ,
										MUX_10_1_IN_2 => UNWINDOWED_443 ,
										MUX_10_1_IN_3 => UNWINDOWED_443 ,
										MUX_10_1_IN_4 => UNWINDOWED_443 ,
										MUX_10_1_IN_5 => UNWINDOWED_443 ,
										MUX_10_1_IN_6 => UNWINDOWED_506 ,
										MUX_10_1_IN_7 => UNWINDOWED_379 ,
										MUX_10_1_IN_8 => UNWINDOWED_379 ,
										MUX_10_1_IN_9 => UNWINDOWED_890 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_445
									);
MUX_REORD_UNIT_446 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_446 ,
										MUX_10_1_IN_1 => UNWINDOWED_445 ,
										MUX_10_1_IN_2 => UNWINDOWED_445 ,
										MUX_10_1_IN_3 => UNWINDOWED_445 ,
										MUX_10_1_IN_4 => UNWINDOWED_445 ,
										MUX_10_1_IN_5 => UNWINDOWED_445 ,
										MUX_10_1_IN_6 => UNWINDOWED_508 ,
										MUX_10_1_IN_7 => UNWINDOWED_381 ,
										MUX_10_1_IN_8 => UNWINDOWED_381 ,
										MUX_10_1_IN_9 => UNWINDOWED_892 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_446
									);
MUX_REORD_UNIT_447 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_447 ,
										MUX_10_1_IN_1 => UNWINDOWED_447 ,
										MUX_10_1_IN_2 => UNWINDOWED_447 ,
										MUX_10_1_IN_3 => UNWINDOWED_447 ,
										MUX_10_1_IN_4 => UNWINDOWED_447 ,
										MUX_10_1_IN_5 => UNWINDOWED_447 ,
										MUX_10_1_IN_6 => UNWINDOWED_510 ,
										MUX_10_1_IN_7 => UNWINDOWED_383 ,
										MUX_10_1_IN_8 => UNWINDOWED_383 ,
										MUX_10_1_IN_9 => UNWINDOWED_894 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_447
									);
MUX_REORD_UNIT_448 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_448 ,
										MUX_10_1_IN_1 => UNWINDOWED_448 ,
										MUX_10_1_IN_2 => UNWINDOWED_448 ,
										MUX_10_1_IN_3 => UNWINDOWED_448 ,
										MUX_10_1_IN_4 => UNWINDOWED_448 ,
										MUX_10_1_IN_5 => UNWINDOWED_448 ,
										MUX_10_1_IN_6 => UNWINDOWED_385 ,
										MUX_10_1_IN_7 => UNWINDOWED_385 ,
										MUX_10_1_IN_8 => UNWINDOWED_385 ,
										MUX_10_1_IN_9 => UNWINDOWED_896 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_448
									);
MUX_REORD_UNIT_449 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_449 ,
										MUX_10_1_IN_1 => UNWINDOWED_450 ,
										MUX_10_1_IN_2 => UNWINDOWED_450 ,
										MUX_10_1_IN_3 => UNWINDOWED_450 ,
										MUX_10_1_IN_4 => UNWINDOWED_450 ,
										MUX_10_1_IN_5 => UNWINDOWED_450 ,
										MUX_10_1_IN_6 => UNWINDOWED_387 ,
										MUX_10_1_IN_7 => UNWINDOWED_387 ,
										MUX_10_1_IN_8 => UNWINDOWED_387 ,
										MUX_10_1_IN_9 => UNWINDOWED_898 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_449
									);
MUX_REORD_UNIT_450 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_450 ,
										MUX_10_1_IN_1 => UNWINDOWED_449 ,
										MUX_10_1_IN_2 => UNWINDOWED_452 ,
										MUX_10_1_IN_3 => UNWINDOWED_452 ,
										MUX_10_1_IN_4 => UNWINDOWED_452 ,
										MUX_10_1_IN_5 => UNWINDOWED_452 ,
										MUX_10_1_IN_6 => UNWINDOWED_389 ,
										MUX_10_1_IN_7 => UNWINDOWED_389 ,
										MUX_10_1_IN_8 => UNWINDOWED_389 ,
										MUX_10_1_IN_9 => UNWINDOWED_900 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_450
									);
MUX_REORD_UNIT_451 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_451 ,
										MUX_10_1_IN_1 => UNWINDOWED_451 ,
										MUX_10_1_IN_2 => UNWINDOWED_454 ,
										MUX_10_1_IN_3 => UNWINDOWED_454 ,
										MUX_10_1_IN_4 => UNWINDOWED_454 ,
										MUX_10_1_IN_5 => UNWINDOWED_454 ,
										MUX_10_1_IN_6 => UNWINDOWED_391 ,
										MUX_10_1_IN_7 => UNWINDOWED_391 ,
										MUX_10_1_IN_8 => UNWINDOWED_391 ,
										MUX_10_1_IN_9 => UNWINDOWED_902 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_451
									);
MUX_REORD_UNIT_452 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_452 ,
										MUX_10_1_IN_1 => UNWINDOWED_452 ,
										MUX_10_1_IN_2 => UNWINDOWED_449 ,
										MUX_10_1_IN_3 => UNWINDOWED_456 ,
										MUX_10_1_IN_4 => UNWINDOWED_456 ,
										MUX_10_1_IN_5 => UNWINDOWED_456 ,
										MUX_10_1_IN_6 => UNWINDOWED_393 ,
										MUX_10_1_IN_7 => UNWINDOWED_393 ,
										MUX_10_1_IN_8 => UNWINDOWED_393 ,
										MUX_10_1_IN_9 => UNWINDOWED_904 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_452
									);
MUX_REORD_UNIT_453 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_453 ,
										MUX_10_1_IN_1 => UNWINDOWED_454 ,
										MUX_10_1_IN_2 => UNWINDOWED_451 ,
										MUX_10_1_IN_3 => UNWINDOWED_458 ,
										MUX_10_1_IN_4 => UNWINDOWED_458 ,
										MUX_10_1_IN_5 => UNWINDOWED_458 ,
										MUX_10_1_IN_6 => UNWINDOWED_395 ,
										MUX_10_1_IN_7 => UNWINDOWED_395 ,
										MUX_10_1_IN_8 => UNWINDOWED_395 ,
										MUX_10_1_IN_9 => UNWINDOWED_906 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_453
									);
MUX_REORD_UNIT_454 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_454 ,
										MUX_10_1_IN_1 => UNWINDOWED_453 ,
										MUX_10_1_IN_2 => UNWINDOWED_453 ,
										MUX_10_1_IN_3 => UNWINDOWED_460 ,
										MUX_10_1_IN_4 => UNWINDOWED_460 ,
										MUX_10_1_IN_5 => UNWINDOWED_460 ,
										MUX_10_1_IN_6 => UNWINDOWED_397 ,
										MUX_10_1_IN_7 => UNWINDOWED_397 ,
										MUX_10_1_IN_8 => UNWINDOWED_397 ,
										MUX_10_1_IN_9 => UNWINDOWED_908 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_454
									);
MUX_REORD_UNIT_455 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_455 ,
										MUX_10_1_IN_1 => UNWINDOWED_455 ,
										MUX_10_1_IN_2 => UNWINDOWED_455 ,
										MUX_10_1_IN_3 => UNWINDOWED_462 ,
										MUX_10_1_IN_4 => UNWINDOWED_462 ,
										MUX_10_1_IN_5 => UNWINDOWED_462 ,
										MUX_10_1_IN_6 => UNWINDOWED_399 ,
										MUX_10_1_IN_7 => UNWINDOWED_399 ,
										MUX_10_1_IN_8 => UNWINDOWED_399 ,
										MUX_10_1_IN_9 => UNWINDOWED_910 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_455
									);
MUX_REORD_UNIT_456 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_456 ,
										MUX_10_1_IN_1 => UNWINDOWED_456 ,
										MUX_10_1_IN_2 => UNWINDOWED_456 ,
										MUX_10_1_IN_3 => UNWINDOWED_449 ,
										MUX_10_1_IN_4 => UNWINDOWED_464 ,
										MUX_10_1_IN_5 => UNWINDOWED_464 ,
										MUX_10_1_IN_6 => UNWINDOWED_401 ,
										MUX_10_1_IN_7 => UNWINDOWED_401 ,
										MUX_10_1_IN_8 => UNWINDOWED_401 ,
										MUX_10_1_IN_9 => UNWINDOWED_912 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_456
									);
MUX_REORD_UNIT_457 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_457 ,
										MUX_10_1_IN_1 => UNWINDOWED_458 ,
										MUX_10_1_IN_2 => UNWINDOWED_458 ,
										MUX_10_1_IN_3 => UNWINDOWED_451 ,
										MUX_10_1_IN_4 => UNWINDOWED_466 ,
										MUX_10_1_IN_5 => UNWINDOWED_466 ,
										MUX_10_1_IN_6 => UNWINDOWED_403 ,
										MUX_10_1_IN_7 => UNWINDOWED_403 ,
										MUX_10_1_IN_8 => UNWINDOWED_403 ,
										MUX_10_1_IN_9 => UNWINDOWED_914 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_457
									);
MUX_REORD_UNIT_458 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_458 ,
										MUX_10_1_IN_1 => UNWINDOWED_457 ,
										MUX_10_1_IN_2 => UNWINDOWED_460 ,
										MUX_10_1_IN_3 => UNWINDOWED_453 ,
										MUX_10_1_IN_4 => UNWINDOWED_468 ,
										MUX_10_1_IN_5 => UNWINDOWED_468 ,
										MUX_10_1_IN_6 => UNWINDOWED_405 ,
										MUX_10_1_IN_7 => UNWINDOWED_405 ,
										MUX_10_1_IN_8 => UNWINDOWED_405 ,
										MUX_10_1_IN_9 => UNWINDOWED_916 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_458
									);
MUX_REORD_UNIT_459 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_459 ,
										MUX_10_1_IN_1 => UNWINDOWED_459 ,
										MUX_10_1_IN_2 => UNWINDOWED_462 ,
										MUX_10_1_IN_3 => UNWINDOWED_455 ,
										MUX_10_1_IN_4 => UNWINDOWED_470 ,
										MUX_10_1_IN_5 => UNWINDOWED_470 ,
										MUX_10_1_IN_6 => UNWINDOWED_407 ,
										MUX_10_1_IN_7 => UNWINDOWED_407 ,
										MUX_10_1_IN_8 => UNWINDOWED_407 ,
										MUX_10_1_IN_9 => UNWINDOWED_918 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_459
									);
MUX_REORD_UNIT_460 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_460 ,
										MUX_10_1_IN_1 => UNWINDOWED_460 ,
										MUX_10_1_IN_2 => UNWINDOWED_457 ,
										MUX_10_1_IN_3 => UNWINDOWED_457 ,
										MUX_10_1_IN_4 => UNWINDOWED_472 ,
										MUX_10_1_IN_5 => UNWINDOWED_472 ,
										MUX_10_1_IN_6 => UNWINDOWED_409 ,
										MUX_10_1_IN_7 => UNWINDOWED_409 ,
										MUX_10_1_IN_8 => UNWINDOWED_409 ,
										MUX_10_1_IN_9 => UNWINDOWED_920 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_460
									);
MUX_REORD_UNIT_461 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_461 ,
										MUX_10_1_IN_1 => UNWINDOWED_462 ,
										MUX_10_1_IN_2 => UNWINDOWED_459 ,
										MUX_10_1_IN_3 => UNWINDOWED_459 ,
										MUX_10_1_IN_4 => UNWINDOWED_474 ,
										MUX_10_1_IN_5 => UNWINDOWED_474 ,
										MUX_10_1_IN_6 => UNWINDOWED_411 ,
										MUX_10_1_IN_7 => UNWINDOWED_411 ,
										MUX_10_1_IN_8 => UNWINDOWED_411 ,
										MUX_10_1_IN_9 => UNWINDOWED_922 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_461
									);
MUX_REORD_UNIT_462 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_462 ,
										MUX_10_1_IN_1 => UNWINDOWED_461 ,
										MUX_10_1_IN_2 => UNWINDOWED_461 ,
										MUX_10_1_IN_3 => UNWINDOWED_461 ,
										MUX_10_1_IN_4 => UNWINDOWED_476 ,
										MUX_10_1_IN_5 => UNWINDOWED_476 ,
										MUX_10_1_IN_6 => UNWINDOWED_413 ,
										MUX_10_1_IN_7 => UNWINDOWED_413 ,
										MUX_10_1_IN_8 => UNWINDOWED_413 ,
										MUX_10_1_IN_9 => UNWINDOWED_924 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_462
									);
MUX_REORD_UNIT_463 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_463 ,
										MUX_10_1_IN_1 => UNWINDOWED_463 ,
										MUX_10_1_IN_2 => UNWINDOWED_463 ,
										MUX_10_1_IN_3 => UNWINDOWED_463 ,
										MUX_10_1_IN_4 => UNWINDOWED_478 ,
										MUX_10_1_IN_5 => UNWINDOWED_478 ,
										MUX_10_1_IN_6 => UNWINDOWED_415 ,
										MUX_10_1_IN_7 => UNWINDOWED_415 ,
										MUX_10_1_IN_8 => UNWINDOWED_415 ,
										MUX_10_1_IN_9 => UNWINDOWED_926 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_463
									);
MUX_REORD_UNIT_464 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_464 ,
										MUX_10_1_IN_1 => UNWINDOWED_464 ,
										MUX_10_1_IN_2 => UNWINDOWED_464 ,
										MUX_10_1_IN_3 => UNWINDOWED_464 ,
										MUX_10_1_IN_4 => UNWINDOWED_449 ,
										MUX_10_1_IN_5 => UNWINDOWED_480 ,
										MUX_10_1_IN_6 => UNWINDOWED_417 ,
										MUX_10_1_IN_7 => UNWINDOWED_417 ,
										MUX_10_1_IN_8 => UNWINDOWED_417 ,
										MUX_10_1_IN_9 => UNWINDOWED_928 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_464
									);
MUX_REORD_UNIT_465 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_465 ,
										MUX_10_1_IN_1 => UNWINDOWED_466 ,
										MUX_10_1_IN_2 => UNWINDOWED_466 ,
										MUX_10_1_IN_3 => UNWINDOWED_466 ,
										MUX_10_1_IN_4 => UNWINDOWED_451 ,
										MUX_10_1_IN_5 => UNWINDOWED_482 ,
										MUX_10_1_IN_6 => UNWINDOWED_419 ,
										MUX_10_1_IN_7 => UNWINDOWED_419 ,
										MUX_10_1_IN_8 => UNWINDOWED_419 ,
										MUX_10_1_IN_9 => UNWINDOWED_930 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_465
									);
MUX_REORD_UNIT_466 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_466 ,
										MUX_10_1_IN_1 => UNWINDOWED_465 ,
										MUX_10_1_IN_2 => UNWINDOWED_468 ,
										MUX_10_1_IN_3 => UNWINDOWED_468 ,
										MUX_10_1_IN_4 => UNWINDOWED_453 ,
										MUX_10_1_IN_5 => UNWINDOWED_484 ,
										MUX_10_1_IN_6 => UNWINDOWED_421 ,
										MUX_10_1_IN_7 => UNWINDOWED_421 ,
										MUX_10_1_IN_8 => UNWINDOWED_421 ,
										MUX_10_1_IN_9 => UNWINDOWED_932 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_466
									);
MUX_REORD_UNIT_467 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_467 ,
										MUX_10_1_IN_1 => UNWINDOWED_467 ,
										MUX_10_1_IN_2 => UNWINDOWED_470 ,
										MUX_10_1_IN_3 => UNWINDOWED_470 ,
										MUX_10_1_IN_4 => UNWINDOWED_455 ,
										MUX_10_1_IN_5 => UNWINDOWED_486 ,
										MUX_10_1_IN_6 => UNWINDOWED_423 ,
										MUX_10_1_IN_7 => UNWINDOWED_423 ,
										MUX_10_1_IN_8 => UNWINDOWED_423 ,
										MUX_10_1_IN_9 => UNWINDOWED_934 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_467
									);
MUX_REORD_UNIT_468 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_468 ,
										MUX_10_1_IN_1 => UNWINDOWED_468 ,
										MUX_10_1_IN_2 => UNWINDOWED_465 ,
										MUX_10_1_IN_3 => UNWINDOWED_472 ,
										MUX_10_1_IN_4 => UNWINDOWED_457 ,
										MUX_10_1_IN_5 => UNWINDOWED_488 ,
										MUX_10_1_IN_6 => UNWINDOWED_425 ,
										MUX_10_1_IN_7 => UNWINDOWED_425 ,
										MUX_10_1_IN_8 => UNWINDOWED_425 ,
										MUX_10_1_IN_9 => UNWINDOWED_936 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_468
									);
MUX_REORD_UNIT_469 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_469 ,
										MUX_10_1_IN_1 => UNWINDOWED_470 ,
										MUX_10_1_IN_2 => UNWINDOWED_467 ,
										MUX_10_1_IN_3 => UNWINDOWED_474 ,
										MUX_10_1_IN_4 => UNWINDOWED_459 ,
										MUX_10_1_IN_5 => UNWINDOWED_490 ,
										MUX_10_1_IN_6 => UNWINDOWED_427 ,
										MUX_10_1_IN_7 => UNWINDOWED_427 ,
										MUX_10_1_IN_8 => UNWINDOWED_427 ,
										MUX_10_1_IN_9 => UNWINDOWED_938 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_469
									);
MUX_REORD_UNIT_470 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_470 ,
										MUX_10_1_IN_1 => UNWINDOWED_469 ,
										MUX_10_1_IN_2 => UNWINDOWED_469 ,
										MUX_10_1_IN_3 => UNWINDOWED_476 ,
										MUX_10_1_IN_4 => UNWINDOWED_461 ,
										MUX_10_1_IN_5 => UNWINDOWED_492 ,
										MUX_10_1_IN_6 => UNWINDOWED_429 ,
										MUX_10_1_IN_7 => UNWINDOWED_429 ,
										MUX_10_1_IN_8 => UNWINDOWED_429 ,
										MUX_10_1_IN_9 => UNWINDOWED_940 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_470
									);
MUX_REORD_UNIT_471 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_471 ,
										MUX_10_1_IN_1 => UNWINDOWED_471 ,
										MUX_10_1_IN_2 => UNWINDOWED_471 ,
										MUX_10_1_IN_3 => UNWINDOWED_478 ,
										MUX_10_1_IN_4 => UNWINDOWED_463 ,
										MUX_10_1_IN_5 => UNWINDOWED_494 ,
										MUX_10_1_IN_6 => UNWINDOWED_431 ,
										MUX_10_1_IN_7 => UNWINDOWED_431 ,
										MUX_10_1_IN_8 => UNWINDOWED_431 ,
										MUX_10_1_IN_9 => UNWINDOWED_942 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_471
									);
MUX_REORD_UNIT_472 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_472 ,
										MUX_10_1_IN_1 => UNWINDOWED_472 ,
										MUX_10_1_IN_2 => UNWINDOWED_472 ,
										MUX_10_1_IN_3 => UNWINDOWED_465 ,
										MUX_10_1_IN_4 => UNWINDOWED_465 ,
										MUX_10_1_IN_5 => UNWINDOWED_496 ,
										MUX_10_1_IN_6 => UNWINDOWED_433 ,
										MUX_10_1_IN_7 => UNWINDOWED_433 ,
										MUX_10_1_IN_8 => UNWINDOWED_433 ,
										MUX_10_1_IN_9 => UNWINDOWED_944 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_472
									);
MUX_REORD_UNIT_473 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_473 ,
										MUX_10_1_IN_1 => UNWINDOWED_474 ,
										MUX_10_1_IN_2 => UNWINDOWED_474 ,
										MUX_10_1_IN_3 => UNWINDOWED_467 ,
										MUX_10_1_IN_4 => UNWINDOWED_467 ,
										MUX_10_1_IN_5 => UNWINDOWED_498 ,
										MUX_10_1_IN_6 => UNWINDOWED_435 ,
										MUX_10_1_IN_7 => UNWINDOWED_435 ,
										MUX_10_1_IN_8 => UNWINDOWED_435 ,
										MUX_10_1_IN_9 => UNWINDOWED_946 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_473
									);
MUX_REORD_UNIT_474 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_474 ,
										MUX_10_1_IN_1 => UNWINDOWED_473 ,
										MUX_10_1_IN_2 => UNWINDOWED_476 ,
										MUX_10_1_IN_3 => UNWINDOWED_469 ,
										MUX_10_1_IN_4 => UNWINDOWED_469 ,
										MUX_10_1_IN_5 => UNWINDOWED_500 ,
										MUX_10_1_IN_6 => UNWINDOWED_437 ,
										MUX_10_1_IN_7 => UNWINDOWED_437 ,
										MUX_10_1_IN_8 => UNWINDOWED_437 ,
										MUX_10_1_IN_9 => UNWINDOWED_948 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_474
									);
MUX_REORD_UNIT_475 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_475 ,
										MUX_10_1_IN_1 => UNWINDOWED_475 ,
										MUX_10_1_IN_2 => UNWINDOWED_478 ,
										MUX_10_1_IN_3 => UNWINDOWED_471 ,
										MUX_10_1_IN_4 => UNWINDOWED_471 ,
										MUX_10_1_IN_5 => UNWINDOWED_502 ,
										MUX_10_1_IN_6 => UNWINDOWED_439 ,
										MUX_10_1_IN_7 => UNWINDOWED_439 ,
										MUX_10_1_IN_8 => UNWINDOWED_439 ,
										MUX_10_1_IN_9 => UNWINDOWED_950 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_475
									);
MUX_REORD_UNIT_476 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_476 ,
										MUX_10_1_IN_1 => UNWINDOWED_476 ,
										MUX_10_1_IN_2 => UNWINDOWED_473 ,
										MUX_10_1_IN_3 => UNWINDOWED_473 ,
										MUX_10_1_IN_4 => UNWINDOWED_473 ,
										MUX_10_1_IN_5 => UNWINDOWED_504 ,
										MUX_10_1_IN_6 => UNWINDOWED_441 ,
										MUX_10_1_IN_7 => UNWINDOWED_441 ,
										MUX_10_1_IN_8 => UNWINDOWED_441 ,
										MUX_10_1_IN_9 => UNWINDOWED_952 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_476
									);
MUX_REORD_UNIT_477 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_477 ,
										MUX_10_1_IN_1 => UNWINDOWED_478 ,
										MUX_10_1_IN_2 => UNWINDOWED_475 ,
										MUX_10_1_IN_3 => UNWINDOWED_475 ,
										MUX_10_1_IN_4 => UNWINDOWED_475 ,
										MUX_10_1_IN_5 => UNWINDOWED_506 ,
										MUX_10_1_IN_6 => UNWINDOWED_443 ,
										MUX_10_1_IN_7 => UNWINDOWED_443 ,
										MUX_10_1_IN_8 => UNWINDOWED_443 ,
										MUX_10_1_IN_9 => UNWINDOWED_954 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_477
									);
MUX_REORD_UNIT_478 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_478 ,
										MUX_10_1_IN_1 => UNWINDOWED_477 ,
										MUX_10_1_IN_2 => UNWINDOWED_477 ,
										MUX_10_1_IN_3 => UNWINDOWED_477 ,
										MUX_10_1_IN_4 => UNWINDOWED_477 ,
										MUX_10_1_IN_5 => UNWINDOWED_508 ,
										MUX_10_1_IN_6 => UNWINDOWED_445 ,
										MUX_10_1_IN_7 => UNWINDOWED_445 ,
										MUX_10_1_IN_8 => UNWINDOWED_445 ,
										MUX_10_1_IN_9 => UNWINDOWED_956 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_478
									);
MUX_REORD_UNIT_479 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_479 ,
										MUX_10_1_IN_1 => UNWINDOWED_479 ,
										MUX_10_1_IN_2 => UNWINDOWED_479 ,
										MUX_10_1_IN_3 => UNWINDOWED_479 ,
										MUX_10_1_IN_4 => UNWINDOWED_479 ,
										MUX_10_1_IN_5 => UNWINDOWED_510 ,
										MUX_10_1_IN_6 => UNWINDOWED_447 ,
										MUX_10_1_IN_7 => UNWINDOWED_447 ,
										MUX_10_1_IN_8 => UNWINDOWED_447 ,
										MUX_10_1_IN_9 => UNWINDOWED_958 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_479
									);
MUX_REORD_UNIT_480 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_480 ,
										MUX_10_1_IN_1 => UNWINDOWED_480 ,
										MUX_10_1_IN_2 => UNWINDOWED_480 ,
										MUX_10_1_IN_3 => UNWINDOWED_480 ,
										MUX_10_1_IN_4 => UNWINDOWED_480 ,
										MUX_10_1_IN_5 => UNWINDOWED_449 ,
										MUX_10_1_IN_6 => UNWINDOWED_449 ,
										MUX_10_1_IN_7 => UNWINDOWED_449 ,
										MUX_10_1_IN_8 => UNWINDOWED_449 ,
										MUX_10_1_IN_9 => UNWINDOWED_960 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_480
									);
MUX_REORD_UNIT_481 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_481 ,
										MUX_10_1_IN_1 => UNWINDOWED_482 ,
										MUX_10_1_IN_2 => UNWINDOWED_482 ,
										MUX_10_1_IN_3 => UNWINDOWED_482 ,
										MUX_10_1_IN_4 => UNWINDOWED_482 ,
										MUX_10_1_IN_5 => UNWINDOWED_451 ,
										MUX_10_1_IN_6 => UNWINDOWED_451 ,
										MUX_10_1_IN_7 => UNWINDOWED_451 ,
										MUX_10_1_IN_8 => UNWINDOWED_451 ,
										MUX_10_1_IN_9 => UNWINDOWED_962 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_481
									);
MUX_REORD_UNIT_482 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_482 ,
										MUX_10_1_IN_1 => UNWINDOWED_481 ,
										MUX_10_1_IN_2 => UNWINDOWED_484 ,
										MUX_10_1_IN_3 => UNWINDOWED_484 ,
										MUX_10_1_IN_4 => UNWINDOWED_484 ,
										MUX_10_1_IN_5 => UNWINDOWED_453 ,
										MUX_10_1_IN_6 => UNWINDOWED_453 ,
										MUX_10_1_IN_7 => UNWINDOWED_453 ,
										MUX_10_1_IN_8 => UNWINDOWED_453 ,
										MUX_10_1_IN_9 => UNWINDOWED_964 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_482
									);
MUX_REORD_UNIT_483 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_483 ,
										MUX_10_1_IN_1 => UNWINDOWED_483 ,
										MUX_10_1_IN_2 => UNWINDOWED_486 ,
										MUX_10_1_IN_3 => UNWINDOWED_486 ,
										MUX_10_1_IN_4 => UNWINDOWED_486 ,
										MUX_10_1_IN_5 => UNWINDOWED_455 ,
										MUX_10_1_IN_6 => UNWINDOWED_455 ,
										MUX_10_1_IN_7 => UNWINDOWED_455 ,
										MUX_10_1_IN_8 => UNWINDOWED_455 ,
										MUX_10_1_IN_9 => UNWINDOWED_966 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_483
									);
MUX_REORD_UNIT_484 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_484 ,
										MUX_10_1_IN_1 => UNWINDOWED_484 ,
										MUX_10_1_IN_2 => UNWINDOWED_481 ,
										MUX_10_1_IN_3 => UNWINDOWED_488 ,
										MUX_10_1_IN_4 => UNWINDOWED_488 ,
										MUX_10_1_IN_5 => UNWINDOWED_457 ,
										MUX_10_1_IN_6 => UNWINDOWED_457 ,
										MUX_10_1_IN_7 => UNWINDOWED_457 ,
										MUX_10_1_IN_8 => UNWINDOWED_457 ,
										MUX_10_1_IN_9 => UNWINDOWED_968 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_484
									);
MUX_REORD_UNIT_485 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_485 ,
										MUX_10_1_IN_1 => UNWINDOWED_486 ,
										MUX_10_1_IN_2 => UNWINDOWED_483 ,
										MUX_10_1_IN_3 => UNWINDOWED_490 ,
										MUX_10_1_IN_4 => UNWINDOWED_490 ,
										MUX_10_1_IN_5 => UNWINDOWED_459 ,
										MUX_10_1_IN_6 => UNWINDOWED_459 ,
										MUX_10_1_IN_7 => UNWINDOWED_459 ,
										MUX_10_1_IN_8 => UNWINDOWED_459 ,
										MUX_10_1_IN_9 => UNWINDOWED_970 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_485
									);
MUX_REORD_UNIT_486 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_486 ,
										MUX_10_1_IN_1 => UNWINDOWED_485 ,
										MUX_10_1_IN_2 => UNWINDOWED_485 ,
										MUX_10_1_IN_3 => UNWINDOWED_492 ,
										MUX_10_1_IN_4 => UNWINDOWED_492 ,
										MUX_10_1_IN_5 => UNWINDOWED_461 ,
										MUX_10_1_IN_6 => UNWINDOWED_461 ,
										MUX_10_1_IN_7 => UNWINDOWED_461 ,
										MUX_10_1_IN_8 => UNWINDOWED_461 ,
										MUX_10_1_IN_9 => UNWINDOWED_972 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_486
									);
MUX_REORD_UNIT_487 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_487 ,
										MUX_10_1_IN_1 => UNWINDOWED_487 ,
										MUX_10_1_IN_2 => UNWINDOWED_487 ,
										MUX_10_1_IN_3 => UNWINDOWED_494 ,
										MUX_10_1_IN_4 => UNWINDOWED_494 ,
										MUX_10_1_IN_5 => UNWINDOWED_463 ,
										MUX_10_1_IN_6 => UNWINDOWED_463 ,
										MUX_10_1_IN_7 => UNWINDOWED_463 ,
										MUX_10_1_IN_8 => UNWINDOWED_463 ,
										MUX_10_1_IN_9 => UNWINDOWED_974 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_487
									);
MUX_REORD_UNIT_488 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_488 ,
										MUX_10_1_IN_1 => UNWINDOWED_488 ,
										MUX_10_1_IN_2 => UNWINDOWED_488 ,
										MUX_10_1_IN_3 => UNWINDOWED_481 ,
										MUX_10_1_IN_4 => UNWINDOWED_496 ,
										MUX_10_1_IN_5 => UNWINDOWED_465 ,
										MUX_10_1_IN_6 => UNWINDOWED_465 ,
										MUX_10_1_IN_7 => UNWINDOWED_465 ,
										MUX_10_1_IN_8 => UNWINDOWED_465 ,
										MUX_10_1_IN_9 => UNWINDOWED_976 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_488
									);
MUX_REORD_UNIT_489 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_489 ,
										MUX_10_1_IN_1 => UNWINDOWED_490 ,
										MUX_10_1_IN_2 => UNWINDOWED_490 ,
										MUX_10_1_IN_3 => UNWINDOWED_483 ,
										MUX_10_1_IN_4 => UNWINDOWED_498 ,
										MUX_10_1_IN_5 => UNWINDOWED_467 ,
										MUX_10_1_IN_6 => UNWINDOWED_467 ,
										MUX_10_1_IN_7 => UNWINDOWED_467 ,
										MUX_10_1_IN_8 => UNWINDOWED_467 ,
										MUX_10_1_IN_9 => UNWINDOWED_978 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_489
									);
MUX_REORD_UNIT_490 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_490 ,
										MUX_10_1_IN_1 => UNWINDOWED_489 ,
										MUX_10_1_IN_2 => UNWINDOWED_492 ,
										MUX_10_1_IN_3 => UNWINDOWED_485 ,
										MUX_10_1_IN_4 => UNWINDOWED_500 ,
										MUX_10_1_IN_5 => UNWINDOWED_469 ,
										MUX_10_1_IN_6 => UNWINDOWED_469 ,
										MUX_10_1_IN_7 => UNWINDOWED_469 ,
										MUX_10_1_IN_8 => UNWINDOWED_469 ,
										MUX_10_1_IN_9 => UNWINDOWED_980 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_490
									);
MUX_REORD_UNIT_491 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_491 ,
										MUX_10_1_IN_1 => UNWINDOWED_491 ,
										MUX_10_1_IN_2 => UNWINDOWED_494 ,
										MUX_10_1_IN_3 => UNWINDOWED_487 ,
										MUX_10_1_IN_4 => UNWINDOWED_502 ,
										MUX_10_1_IN_5 => UNWINDOWED_471 ,
										MUX_10_1_IN_6 => UNWINDOWED_471 ,
										MUX_10_1_IN_7 => UNWINDOWED_471 ,
										MUX_10_1_IN_8 => UNWINDOWED_471 ,
										MUX_10_1_IN_9 => UNWINDOWED_982 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_491
									);
MUX_REORD_UNIT_492 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_492 ,
										MUX_10_1_IN_1 => UNWINDOWED_492 ,
										MUX_10_1_IN_2 => UNWINDOWED_489 ,
										MUX_10_1_IN_3 => UNWINDOWED_489 ,
										MUX_10_1_IN_4 => UNWINDOWED_504 ,
										MUX_10_1_IN_5 => UNWINDOWED_473 ,
										MUX_10_1_IN_6 => UNWINDOWED_473 ,
										MUX_10_1_IN_7 => UNWINDOWED_473 ,
										MUX_10_1_IN_8 => UNWINDOWED_473 ,
										MUX_10_1_IN_9 => UNWINDOWED_984 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_492
									);
MUX_REORD_UNIT_493 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_493 ,
										MUX_10_1_IN_1 => UNWINDOWED_494 ,
										MUX_10_1_IN_2 => UNWINDOWED_491 ,
										MUX_10_1_IN_3 => UNWINDOWED_491 ,
										MUX_10_1_IN_4 => UNWINDOWED_506 ,
										MUX_10_1_IN_5 => UNWINDOWED_475 ,
										MUX_10_1_IN_6 => UNWINDOWED_475 ,
										MUX_10_1_IN_7 => UNWINDOWED_475 ,
										MUX_10_1_IN_8 => UNWINDOWED_475 ,
										MUX_10_1_IN_9 => UNWINDOWED_986 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_493
									);
MUX_REORD_UNIT_494 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_494 ,
										MUX_10_1_IN_1 => UNWINDOWED_493 ,
										MUX_10_1_IN_2 => UNWINDOWED_493 ,
										MUX_10_1_IN_3 => UNWINDOWED_493 ,
										MUX_10_1_IN_4 => UNWINDOWED_508 ,
										MUX_10_1_IN_5 => UNWINDOWED_477 ,
										MUX_10_1_IN_6 => UNWINDOWED_477 ,
										MUX_10_1_IN_7 => UNWINDOWED_477 ,
										MUX_10_1_IN_8 => UNWINDOWED_477 ,
										MUX_10_1_IN_9 => UNWINDOWED_988 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_494
									);
MUX_REORD_UNIT_495 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_495 ,
										MUX_10_1_IN_1 => UNWINDOWED_495 ,
										MUX_10_1_IN_2 => UNWINDOWED_495 ,
										MUX_10_1_IN_3 => UNWINDOWED_495 ,
										MUX_10_1_IN_4 => UNWINDOWED_510 ,
										MUX_10_1_IN_5 => UNWINDOWED_479 ,
										MUX_10_1_IN_6 => UNWINDOWED_479 ,
										MUX_10_1_IN_7 => UNWINDOWED_479 ,
										MUX_10_1_IN_8 => UNWINDOWED_479 ,
										MUX_10_1_IN_9 => UNWINDOWED_990 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_495
									);
MUX_REORD_UNIT_496 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_496 ,
										MUX_10_1_IN_1 => UNWINDOWED_496 ,
										MUX_10_1_IN_2 => UNWINDOWED_496 ,
										MUX_10_1_IN_3 => UNWINDOWED_496 ,
										MUX_10_1_IN_4 => UNWINDOWED_481 ,
										MUX_10_1_IN_5 => UNWINDOWED_481 ,
										MUX_10_1_IN_6 => UNWINDOWED_481 ,
										MUX_10_1_IN_7 => UNWINDOWED_481 ,
										MUX_10_1_IN_8 => UNWINDOWED_481 ,
										MUX_10_1_IN_9 => UNWINDOWED_992 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_496
									);
MUX_REORD_UNIT_497 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_497 ,
										MUX_10_1_IN_1 => UNWINDOWED_498 ,
										MUX_10_1_IN_2 => UNWINDOWED_498 ,
										MUX_10_1_IN_3 => UNWINDOWED_498 ,
										MUX_10_1_IN_4 => UNWINDOWED_483 ,
										MUX_10_1_IN_5 => UNWINDOWED_483 ,
										MUX_10_1_IN_6 => UNWINDOWED_483 ,
										MUX_10_1_IN_7 => UNWINDOWED_483 ,
										MUX_10_1_IN_8 => UNWINDOWED_483 ,
										MUX_10_1_IN_9 => UNWINDOWED_994 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_497
									);
MUX_REORD_UNIT_498 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_498 ,
										MUX_10_1_IN_1 => UNWINDOWED_497 ,
										MUX_10_1_IN_2 => UNWINDOWED_500 ,
										MUX_10_1_IN_3 => UNWINDOWED_500 ,
										MUX_10_1_IN_4 => UNWINDOWED_485 ,
										MUX_10_1_IN_5 => UNWINDOWED_485 ,
										MUX_10_1_IN_6 => UNWINDOWED_485 ,
										MUX_10_1_IN_7 => UNWINDOWED_485 ,
										MUX_10_1_IN_8 => UNWINDOWED_485 ,
										MUX_10_1_IN_9 => UNWINDOWED_996 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_498
									);
MUX_REORD_UNIT_499 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_499 ,
										MUX_10_1_IN_1 => UNWINDOWED_499 ,
										MUX_10_1_IN_2 => UNWINDOWED_502 ,
										MUX_10_1_IN_3 => UNWINDOWED_502 ,
										MUX_10_1_IN_4 => UNWINDOWED_487 ,
										MUX_10_1_IN_5 => UNWINDOWED_487 ,
										MUX_10_1_IN_6 => UNWINDOWED_487 ,
										MUX_10_1_IN_7 => UNWINDOWED_487 ,
										MUX_10_1_IN_8 => UNWINDOWED_487 ,
										MUX_10_1_IN_9 => UNWINDOWED_998 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_499
									);
MUX_REORD_UNIT_500 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_500 ,
										MUX_10_1_IN_1 => UNWINDOWED_500 ,
										MUX_10_1_IN_2 => UNWINDOWED_497 ,
										MUX_10_1_IN_3 => UNWINDOWED_504 ,
										MUX_10_1_IN_4 => UNWINDOWED_489 ,
										MUX_10_1_IN_5 => UNWINDOWED_489 ,
										MUX_10_1_IN_6 => UNWINDOWED_489 ,
										MUX_10_1_IN_7 => UNWINDOWED_489 ,
										MUX_10_1_IN_8 => UNWINDOWED_489 ,
										MUX_10_1_IN_9 => UNWINDOWED_1000 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_500
									);
MUX_REORD_UNIT_501 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_501 ,
										MUX_10_1_IN_1 => UNWINDOWED_502 ,
										MUX_10_1_IN_2 => UNWINDOWED_499 ,
										MUX_10_1_IN_3 => UNWINDOWED_506 ,
										MUX_10_1_IN_4 => UNWINDOWED_491 ,
										MUX_10_1_IN_5 => UNWINDOWED_491 ,
										MUX_10_1_IN_6 => UNWINDOWED_491 ,
										MUX_10_1_IN_7 => UNWINDOWED_491 ,
										MUX_10_1_IN_8 => UNWINDOWED_491 ,
										MUX_10_1_IN_9 => UNWINDOWED_1002 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_501
									);
MUX_REORD_UNIT_502 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_502 ,
										MUX_10_1_IN_1 => UNWINDOWED_501 ,
										MUX_10_1_IN_2 => UNWINDOWED_501 ,
										MUX_10_1_IN_3 => UNWINDOWED_508 ,
										MUX_10_1_IN_4 => UNWINDOWED_493 ,
										MUX_10_1_IN_5 => UNWINDOWED_493 ,
										MUX_10_1_IN_6 => UNWINDOWED_493 ,
										MUX_10_1_IN_7 => UNWINDOWED_493 ,
										MUX_10_1_IN_8 => UNWINDOWED_493 ,
										MUX_10_1_IN_9 => UNWINDOWED_1004 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_502
									);
MUX_REORD_UNIT_503 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_503 ,
										MUX_10_1_IN_1 => UNWINDOWED_503 ,
										MUX_10_1_IN_2 => UNWINDOWED_503 ,
										MUX_10_1_IN_3 => UNWINDOWED_510 ,
										MUX_10_1_IN_4 => UNWINDOWED_495 ,
										MUX_10_1_IN_5 => UNWINDOWED_495 ,
										MUX_10_1_IN_6 => UNWINDOWED_495 ,
										MUX_10_1_IN_7 => UNWINDOWED_495 ,
										MUX_10_1_IN_8 => UNWINDOWED_495 ,
										MUX_10_1_IN_9 => UNWINDOWED_1006 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_503
									);
MUX_REORD_UNIT_504 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_504 ,
										MUX_10_1_IN_1 => UNWINDOWED_504 ,
										MUX_10_1_IN_2 => UNWINDOWED_504 ,
										MUX_10_1_IN_3 => UNWINDOWED_497 ,
										MUX_10_1_IN_4 => UNWINDOWED_497 ,
										MUX_10_1_IN_5 => UNWINDOWED_497 ,
										MUX_10_1_IN_6 => UNWINDOWED_497 ,
										MUX_10_1_IN_7 => UNWINDOWED_497 ,
										MUX_10_1_IN_8 => UNWINDOWED_497 ,
										MUX_10_1_IN_9 => UNWINDOWED_1008 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_504
									);
MUX_REORD_UNIT_505 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_505 ,
										MUX_10_1_IN_1 => UNWINDOWED_506 ,
										MUX_10_1_IN_2 => UNWINDOWED_506 ,
										MUX_10_1_IN_3 => UNWINDOWED_499 ,
										MUX_10_1_IN_4 => UNWINDOWED_499 ,
										MUX_10_1_IN_5 => UNWINDOWED_499 ,
										MUX_10_1_IN_6 => UNWINDOWED_499 ,
										MUX_10_1_IN_7 => UNWINDOWED_499 ,
										MUX_10_1_IN_8 => UNWINDOWED_499 ,
										MUX_10_1_IN_9 => UNWINDOWED_1010 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_505
									);
MUX_REORD_UNIT_506 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_506 ,
										MUX_10_1_IN_1 => UNWINDOWED_505 ,
										MUX_10_1_IN_2 => UNWINDOWED_508 ,
										MUX_10_1_IN_3 => UNWINDOWED_501 ,
										MUX_10_1_IN_4 => UNWINDOWED_501 ,
										MUX_10_1_IN_5 => UNWINDOWED_501 ,
										MUX_10_1_IN_6 => UNWINDOWED_501 ,
										MUX_10_1_IN_7 => UNWINDOWED_501 ,
										MUX_10_1_IN_8 => UNWINDOWED_501 ,
										MUX_10_1_IN_9 => UNWINDOWED_1012 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_506
									);
MUX_REORD_UNIT_507 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_507 ,
										MUX_10_1_IN_1 => UNWINDOWED_507 ,
										MUX_10_1_IN_2 => UNWINDOWED_510 ,
										MUX_10_1_IN_3 => UNWINDOWED_503 ,
										MUX_10_1_IN_4 => UNWINDOWED_503 ,
										MUX_10_1_IN_5 => UNWINDOWED_503 ,
										MUX_10_1_IN_6 => UNWINDOWED_503 ,
										MUX_10_1_IN_7 => UNWINDOWED_503 ,
										MUX_10_1_IN_8 => UNWINDOWED_503 ,
										MUX_10_1_IN_9 => UNWINDOWED_1014 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_507
									);
MUX_REORD_UNIT_508 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_508 ,
										MUX_10_1_IN_1 => UNWINDOWED_508 ,
										MUX_10_1_IN_2 => UNWINDOWED_505 ,
										MUX_10_1_IN_3 => UNWINDOWED_505 ,
										MUX_10_1_IN_4 => UNWINDOWED_505 ,
										MUX_10_1_IN_5 => UNWINDOWED_505 ,
										MUX_10_1_IN_6 => UNWINDOWED_505 ,
										MUX_10_1_IN_7 => UNWINDOWED_505 ,
										MUX_10_1_IN_8 => UNWINDOWED_505 ,
										MUX_10_1_IN_9 => UNWINDOWED_1016 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_508
									);
MUX_REORD_UNIT_509 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_509 ,
										MUX_10_1_IN_1 => UNWINDOWED_510 ,
										MUX_10_1_IN_2 => UNWINDOWED_507 ,
										MUX_10_1_IN_3 => UNWINDOWED_507 ,
										MUX_10_1_IN_4 => UNWINDOWED_507 ,
										MUX_10_1_IN_5 => UNWINDOWED_507 ,
										MUX_10_1_IN_6 => UNWINDOWED_507 ,
										MUX_10_1_IN_7 => UNWINDOWED_507 ,
										MUX_10_1_IN_8 => UNWINDOWED_507 ,
										MUX_10_1_IN_9 => UNWINDOWED_1018 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_509
									);
MUX_REORD_UNIT_510 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_510 ,
										MUX_10_1_IN_1 => UNWINDOWED_509 ,
										MUX_10_1_IN_2 => UNWINDOWED_509 ,
										MUX_10_1_IN_3 => UNWINDOWED_509 ,
										MUX_10_1_IN_4 => UNWINDOWED_509 ,
										MUX_10_1_IN_5 => UNWINDOWED_509 ,
										MUX_10_1_IN_6 => UNWINDOWED_509 ,
										MUX_10_1_IN_7 => UNWINDOWED_509 ,
										MUX_10_1_IN_8 => UNWINDOWED_509 ,
										MUX_10_1_IN_9 => UNWINDOWED_1020 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_510
									);
MUX_REORD_UNIT_511 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_511 ,
										MUX_10_1_IN_1 => UNWINDOWED_511 ,
										MUX_10_1_IN_2 => UNWINDOWED_511 ,
										MUX_10_1_IN_3 => UNWINDOWED_511 ,
										MUX_10_1_IN_4 => UNWINDOWED_511 ,
										MUX_10_1_IN_5 => UNWINDOWED_511 ,
										MUX_10_1_IN_6 => UNWINDOWED_511 ,
										MUX_10_1_IN_7 => UNWINDOWED_511 ,
										MUX_10_1_IN_8 => UNWINDOWED_511 ,
										MUX_10_1_IN_9 => UNWINDOWED_1022 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_511
									);
MUX_REORD_UNIT_512 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_512 ,
										MUX_10_1_IN_1 => UNWINDOWED_512 ,
										MUX_10_1_IN_2 => UNWINDOWED_512 ,
										MUX_10_1_IN_3 => UNWINDOWED_512 ,
										MUX_10_1_IN_4 => UNWINDOWED_512 ,
										MUX_10_1_IN_5 => UNWINDOWED_512 ,
										MUX_10_1_IN_6 => UNWINDOWED_512 ,
										MUX_10_1_IN_7 => UNWINDOWED_512 ,
										MUX_10_1_IN_8 => UNWINDOWED_512 ,
										MUX_10_1_IN_9 => UNWINDOWED_1 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_512
									);
MUX_REORD_UNIT_513 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_513 ,
										MUX_10_1_IN_1 => UNWINDOWED_514 ,
										MUX_10_1_IN_2 => UNWINDOWED_514 ,
										MUX_10_1_IN_3 => UNWINDOWED_514 ,
										MUX_10_1_IN_4 => UNWINDOWED_514 ,
										MUX_10_1_IN_5 => UNWINDOWED_514 ,
										MUX_10_1_IN_6 => UNWINDOWED_514 ,
										MUX_10_1_IN_7 => UNWINDOWED_514 ,
										MUX_10_1_IN_8 => UNWINDOWED_514 ,
										MUX_10_1_IN_9 => UNWINDOWED_3 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_513
									);
MUX_REORD_UNIT_514 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_514 ,
										MUX_10_1_IN_1 => UNWINDOWED_513 ,
										MUX_10_1_IN_2 => UNWINDOWED_516 ,
										MUX_10_1_IN_3 => UNWINDOWED_516 ,
										MUX_10_1_IN_4 => UNWINDOWED_516 ,
										MUX_10_1_IN_5 => UNWINDOWED_516 ,
										MUX_10_1_IN_6 => UNWINDOWED_516 ,
										MUX_10_1_IN_7 => UNWINDOWED_516 ,
										MUX_10_1_IN_8 => UNWINDOWED_516 ,
										MUX_10_1_IN_9 => UNWINDOWED_5 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_514
									);
MUX_REORD_UNIT_515 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_515 ,
										MUX_10_1_IN_1 => UNWINDOWED_515 ,
										MUX_10_1_IN_2 => UNWINDOWED_518 ,
										MUX_10_1_IN_3 => UNWINDOWED_518 ,
										MUX_10_1_IN_4 => UNWINDOWED_518 ,
										MUX_10_1_IN_5 => UNWINDOWED_518 ,
										MUX_10_1_IN_6 => UNWINDOWED_518 ,
										MUX_10_1_IN_7 => UNWINDOWED_518 ,
										MUX_10_1_IN_8 => UNWINDOWED_518 ,
										MUX_10_1_IN_9 => UNWINDOWED_7 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_515
									);
MUX_REORD_UNIT_516 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_516 ,
										MUX_10_1_IN_1 => UNWINDOWED_516 ,
										MUX_10_1_IN_2 => UNWINDOWED_513 ,
										MUX_10_1_IN_3 => UNWINDOWED_520 ,
										MUX_10_1_IN_4 => UNWINDOWED_520 ,
										MUX_10_1_IN_5 => UNWINDOWED_520 ,
										MUX_10_1_IN_6 => UNWINDOWED_520 ,
										MUX_10_1_IN_7 => UNWINDOWED_520 ,
										MUX_10_1_IN_8 => UNWINDOWED_520 ,
										MUX_10_1_IN_9 => UNWINDOWED_9 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_516
									);
MUX_REORD_UNIT_517 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_517 ,
										MUX_10_1_IN_1 => UNWINDOWED_518 ,
										MUX_10_1_IN_2 => UNWINDOWED_515 ,
										MUX_10_1_IN_3 => UNWINDOWED_522 ,
										MUX_10_1_IN_4 => UNWINDOWED_522 ,
										MUX_10_1_IN_5 => UNWINDOWED_522 ,
										MUX_10_1_IN_6 => UNWINDOWED_522 ,
										MUX_10_1_IN_7 => UNWINDOWED_522 ,
										MUX_10_1_IN_8 => UNWINDOWED_522 ,
										MUX_10_1_IN_9 => UNWINDOWED_11 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_517
									);
MUX_REORD_UNIT_518 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_518 ,
										MUX_10_1_IN_1 => UNWINDOWED_517 ,
										MUX_10_1_IN_2 => UNWINDOWED_517 ,
										MUX_10_1_IN_3 => UNWINDOWED_524 ,
										MUX_10_1_IN_4 => UNWINDOWED_524 ,
										MUX_10_1_IN_5 => UNWINDOWED_524 ,
										MUX_10_1_IN_6 => UNWINDOWED_524 ,
										MUX_10_1_IN_7 => UNWINDOWED_524 ,
										MUX_10_1_IN_8 => UNWINDOWED_524 ,
										MUX_10_1_IN_9 => UNWINDOWED_13 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_518
									);
MUX_REORD_UNIT_519 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_519 ,
										MUX_10_1_IN_1 => UNWINDOWED_519 ,
										MUX_10_1_IN_2 => UNWINDOWED_519 ,
										MUX_10_1_IN_3 => UNWINDOWED_526 ,
										MUX_10_1_IN_4 => UNWINDOWED_526 ,
										MUX_10_1_IN_5 => UNWINDOWED_526 ,
										MUX_10_1_IN_6 => UNWINDOWED_526 ,
										MUX_10_1_IN_7 => UNWINDOWED_526 ,
										MUX_10_1_IN_8 => UNWINDOWED_526 ,
										MUX_10_1_IN_9 => UNWINDOWED_15 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_519
									);
MUX_REORD_UNIT_520 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_520 ,
										MUX_10_1_IN_1 => UNWINDOWED_520 ,
										MUX_10_1_IN_2 => UNWINDOWED_520 ,
										MUX_10_1_IN_3 => UNWINDOWED_513 ,
										MUX_10_1_IN_4 => UNWINDOWED_528 ,
										MUX_10_1_IN_5 => UNWINDOWED_528 ,
										MUX_10_1_IN_6 => UNWINDOWED_528 ,
										MUX_10_1_IN_7 => UNWINDOWED_528 ,
										MUX_10_1_IN_8 => UNWINDOWED_528 ,
										MUX_10_1_IN_9 => UNWINDOWED_17 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_520
									);
MUX_REORD_UNIT_521 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_521 ,
										MUX_10_1_IN_1 => UNWINDOWED_522 ,
										MUX_10_1_IN_2 => UNWINDOWED_522 ,
										MUX_10_1_IN_3 => UNWINDOWED_515 ,
										MUX_10_1_IN_4 => UNWINDOWED_530 ,
										MUX_10_1_IN_5 => UNWINDOWED_530 ,
										MUX_10_1_IN_6 => UNWINDOWED_530 ,
										MUX_10_1_IN_7 => UNWINDOWED_530 ,
										MUX_10_1_IN_8 => UNWINDOWED_530 ,
										MUX_10_1_IN_9 => UNWINDOWED_19 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_521
									);
MUX_REORD_UNIT_522 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_522 ,
										MUX_10_1_IN_1 => UNWINDOWED_521 ,
										MUX_10_1_IN_2 => UNWINDOWED_524 ,
										MUX_10_1_IN_3 => UNWINDOWED_517 ,
										MUX_10_1_IN_4 => UNWINDOWED_532 ,
										MUX_10_1_IN_5 => UNWINDOWED_532 ,
										MUX_10_1_IN_6 => UNWINDOWED_532 ,
										MUX_10_1_IN_7 => UNWINDOWED_532 ,
										MUX_10_1_IN_8 => UNWINDOWED_532 ,
										MUX_10_1_IN_9 => UNWINDOWED_21 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_522
									);
MUX_REORD_UNIT_523 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_523 ,
										MUX_10_1_IN_1 => UNWINDOWED_523 ,
										MUX_10_1_IN_2 => UNWINDOWED_526 ,
										MUX_10_1_IN_3 => UNWINDOWED_519 ,
										MUX_10_1_IN_4 => UNWINDOWED_534 ,
										MUX_10_1_IN_5 => UNWINDOWED_534 ,
										MUX_10_1_IN_6 => UNWINDOWED_534 ,
										MUX_10_1_IN_7 => UNWINDOWED_534 ,
										MUX_10_1_IN_8 => UNWINDOWED_534 ,
										MUX_10_1_IN_9 => UNWINDOWED_23 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_523
									);
MUX_REORD_UNIT_524 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_524 ,
										MUX_10_1_IN_1 => UNWINDOWED_524 ,
										MUX_10_1_IN_2 => UNWINDOWED_521 ,
										MUX_10_1_IN_3 => UNWINDOWED_521 ,
										MUX_10_1_IN_4 => UNWINDOWED_536 ,
										MUX_10_1_IN_5 => UNWINDOWED_536 ,
										MUX_10_1_IN_6 => UNWINDOWED_536 ,
										MUX_10_1_IN_7 => UNWINDOWED_536 ,
										MUX_10_1_IN_8 => UNWINDOWED_536 ,
										MUX_10_1_IN_9 => UNWINDOWED_25 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_524
									);
MUX_REORD_UNIT_525 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_525 ,
										MUX_10_1_IN_1 => UNWINDOWED_526 ,
										MUX_10_1_IN_2 => UNWINDOWED_523 ,
										MUX_10_1_IN_3 => UNWINDOWED_523 ,
										MUX_10_1_IN_4 => UNWINDOWED_538 ,
										MUX_10_1_IN_5 => UNWINDOWED_538 ,
										MUX_10_1_IN_6 => UNWINDOWED_538 ,
										MUX_10_1_IN_7 => UNWINDOWED_538 ,
										MUX_10_1_IN_8 => UNWINDOWED_538 ,
										MUX_10_1_IN_9 => UNWINDOWED_27 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_525
									);
MUX_REORD_UNIT_526 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_526 ,
										MUX_10_1_IN_1 => UNWINDOWED_525 ,
										MUX_10_1_IN_2 => UNWINDOWED_525 ,
										MUX_10_1_IN_3 => UNWINDOWED_525 ,
										MUX_10_1_IN_4 => UNWINDOWED_540 ,
										MUX_10_1_IN_5 => UNWINDOWED_540 ,
										MUX_10_1_IN_6 => UNWINDOWED_540 ,
										MUX_10_1_IN_7 => UNWINDOWED_540 ,
										MUX_10_1_IN_8 => UNWINDOWED_540 ,
										MUX_10_1_IN_9 => UNWINDOWED_29 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_526
									);
MUX_REORD_UNIT_527 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_527 ,
										MUX_10_1_IN_1 => UNWINDOWED_527 ,
										MUX_10_1_IN_2 => UNWINDOWED_527 ,
										MUX_10_1_IN_3 => UNWINDOWED_527 ,
										MUX_10_1_IN_4 => UNWINDOWED_542 ,
										MUX_10_1_IN_5 => UNWINDOWED_542 ,
										MUX_10_1_IN_6 => UNWINDOWED_542 ,
										MUX_10_1_IN_7 => UNWINDOWED_542 ,
										MUX_10_1_IN_8 => UNWINDOWED_542 ,
										MUX_10_1_IN_9 => UNWINDOWED_31 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_527
									);
MUX_REORD_UNIT_528 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_528 ,
										MUX_10_1_IN_1 => UNWINDOWED_528 ,
										MUX_10_1_IN_2 => UNWINDOWED_528 ,
										MUX_10_1_IN_3 => UNWINDOWED_528 ,
										MUX_10_1_IN_4 => UNWINDOWED_513 ,
										MUX_10_1_IN_5 => UNWINDOWED_544 ,
										MUX_10_1_IN_6 => UNWINDOWED_544 ,
										MUX_10_1_IN_7 => UNWINDOWED_544 ,
										MUX_10_1_IN_8 => UNWINDOWED_544 ,
										MUX_10_1_IN_9 => UNWINDOWED_33 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_528
									);
MUX_REORD_UNIT_529 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_529 ,
										MUX_10_1_IN_1 => UNWINDOWED_530 ,
										MUX_10_1_IN_2 => UNWINDOWED_530 ,
										MUX_10_1_IN_3 => UNWINDOWED_530 ,
										MUX_10_1_IN_4 => UNWINDOWED_515 ,
										MUX_10_1_IN_5 => UNWINDOWED_546 ,
										MUX_10_1_IN_6 => UNWINDOWED_546 ,
										MUX_10_1_IN_7 => UNWINDOWED_546 ,
										MUX_10_1_IN_8 => UNWINDOWED_546 ,
										MUX_10_1_IN_9 => UNWINDOWED_35 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_529
									);
MUX_REORD_UNIT_530 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_530 ,
										MUX_10_1_IN_1 => UNWINDOWED_529 ,
										MUX_10_1_IN_2 => UNWINDOWED_532 ,
										MUX_10_1_IN_3 => UNWINDOWED_532 ,
										MUX_10_1_IN_4 => UNWINDOWED_517 ,
										MUX_10_1_IN_5 => UNWINDOWED_548 ,
										MUX_10_1_IN_6 => UNWINDOWED_548 ,
										MUX_10_1_IN_7 => UNWINDOWED_548 ,
										MUX_10_1_IN_8 => UNWINDOWED_548 ,
										MUX_10_1_IN_9 => UNWINDOWED_37 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_530
									);
MUX_REORD_UNIT_531 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_531 ,
										MUX_10_1_IN_1 => UNWINDOWED_531 ,
										MUX_10_1_IN_2 => UNWINDOWED_534 ,
										MUX_10_1_IN_3 => UNWINDOWED_534 ,
										MUX_10_1_IN_4 => UNWINDOWED_519 ,
										MUX_10_1_IN_5 => UNWINDOWED_550 ,
										MUX_10_1_IN_6 => UNWINDOWED_550 ,
										MUX_10_1_IN_7 => UNWINDOWED_550 ,
										MUX_10_1_IN_8 => UNWINDOWED_550 ,
										MUX_10_1_IN_9 => UNWINDOWED_39 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_531
									);
MUX_REORD_UNIT_532 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_532 ,
										MUX_10_1_IN_1 => UNWINDOWED_532 ,
										MUX_10_1_IN_2 => UNWINDOWED_529 ,
										MUX_10_1_IN_3 => UNWINDOWED_536 ,
										MUX_10_1_IN_4 => UNWINDOWED_521 ,
										MUX_10_1_IN_5 => UNWINDOWED_552 ,
										MUX_10_1_IN_6 => UNWINDOWED_552 ,
										MUX_10_1_IN_7 => UNWINDOWED_552 ,
										MUX_10_1_IN_8 => UNWINDOWED_552 ,
										MUX_10_1_IN_9 => UNWINDOWED_41 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_532
									);
MUX_REORD_UNIT_533 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_533 ,
										MUX_10_1_IN_1 => UNWINDOWED_534 ,
										MUX_10_1_IN_2 => UNWINDOWED_531 ,
										MUX_10_1_IN_3 => UNWINDOWED_538 ,
										MUX_10_1_IN_4 => UNWINDOWED_523 ,
										MUX_10_1_IN_5 => UNWINDOWED_554 ,
										MUX_10_1_IN_6 => UNWINDOWED_554 ,
										MUX_10_1_IN_7 => UNWINDOWED_554 ,
										MUX_10_1_IN_8 => UNWINDOWED_554 ,
										MUX_10_1_IN_9 => UNWINDOWED_43 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_533
									);
MUX_REORD_UNIT_534 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_534 ,
										MUX_10_1_IN_1 => UNWINDOWED_533 ,
										MUX_10_1_IN_2 => UNWINDOWED_533 ,
										MUX_10_1_IN_3 => UNWINDOWED_540 ,
										MUX_10_1_IN_4 => UNWINDOWED_525 ,
										MUX_10_1_IN_5 => UNWINDOWED_556 ,
										MUX_10_1_IN_6 => UNWINDOWED_556 ,
										MUX_10_1_IN_7 => UNWINDOWED_556 ,
										MUX_10_1_IN_8 => UNWINDOWED_556 ,
										MUX_10_1_IN_9 => UNWINDOWED_45 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_534
									);
MUX_REORD_UNIT_535 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_535 ,
										MUX_10_1_IN_1 => UNWINDOWED_535 ,
										MUX_10_1_IN_2 => UNWINDOWED_535 ,
										MUX_10_1_IN_3 => UNWINDOWED_542 ,
										MUX_10_1_IN_4 => UNWINDOWED_527 ,
										MUX_10_1_IN_5 => UNWINDOWED_558 ,
										MUX_10_1_IN_6 => UNWINDOWED_558 ,
										MUX_10_1_IN_7 => UNWINDOWED_558 ,
										MUX_10_1_IN_8 => UNWINDOWED_558 ,
										MUX_10_1_IN_9 => UNWINDOWED_47 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_535
									);
MUX_REORD_UNIT_536 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_536 ,
										MUX_10_1_IN_1 => UNWINDOWED_536 ,
										MUX_10_1_IN_2 => UNWINDOWED_536 ,
										MUX_10_1_IN_3 => UNWINDOWED_529 ,
										MUX_10_1_IN_4 => UNWINDOWED_529 ,
										MUX_10_1_IN_5 => UNWINDOWED_560 ,
										MUX_10_1_IN_6 => UNWINDOWED_560 ,
										MUX_10_1_IN_7 => UNWINDOWED_560 ,
										MUX_10_1_IN_8 => UNWINDOWED_560 ,
										MUX_10_1_IN_9 => UNWINDOWED_49 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_536
									);
MUX_REORD_UNIT_537 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_537 ,
										MUX_10_1_IN_1 => UNWINDOWED_538 ,
										MUX_10_1_IN_2 => UNWINDOWED_538 ,
										MUX_10_1_IN_3 => UNWINDOWED_531 ,
										MUX_10_1_IN_4 => UNWINDOWED_531 ,
										MUX_10_1_IN_5 => UNWINDOWED_562 ,
										MUX_10_1_IN_6 => UNWINDOWED_562 ,
										MUX_10_1_IN_7 => UNWINDOWED_562 ,
										MUX_10_1_IN_8 => UNWINDOWED_562 ,
										MUX_10_1_IN_9 => UNWINDOWED_51 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_537
									);
MUX_REORD_UNIT_538 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_538 ,
										MUX_10_1_IN_1 => UNWINDOWED_537 ,
										MUX_10_1_IN_2 => UNWINDOWED_540 ,
										MUX_10_1_IN_3 => UNWINDOWED_533 ,
										MUX_10_1_IN_4 => UNWINDOWED_533 ,
										MUX_10_1_IN_5 => UNWINDOWED_564 ,
										MUX_10_1_IN_6 => UNWINDOWED_564 ,
										MUX_10_1_IN_7 => UNWINDOWED_564 ,
										MUX_10_1_IN_8 => UNWINDOWED_564 ,
										MUX_10_1_IN_9 => UNWINDOWED_53 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_538
									);
MUX_REORD_UNIT_539 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_539 ,
										MUX_10_1_IN_1 => UNWINDOWED_539 ,
										MUX_10_1_IN_2 => UNWINDOWED_542 ,
										MUX_10_1_IN_3 => UNWINDOWED_535 ,
										MUX_10_1_IN_4 => UNWINDOWED_535 ,
										MUX_10_1_IN_5 => UNWINDOWED_566 ,
										MUX_10_1_IN_6 => UNWINDOWED_566 ,
										MUX_10_1_IN_7 => UNWINDOWED_566 ,
										MUX_10_1_IN_8 => UNWINDOWED_566 ,
										MUX_10_1_IN_9 => UNWINDOWED_55 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_539
									);
MUX_REORD_UNIT_540 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_540 ,
										MUX_10_1_IN_1 => UNWINDOWED_540 ,
										MUX_10_1_IN_2 => UNWINDOWED_537 ,
										MUX_10_1_IN_3 => UNWINDOWED_537 ,
										MUX_10_1_IN_4 => UNWINDOWED_537 ,
										MUX_10_1_IN_5 => UNWINDOWED_568 ,
										MUX_10_1_IN_6 => UNWINDOWED_568 ,
										MUX_10_1_IN_7 => UNWINDOWED_568 ,
										MUX_10_1_IN_8 => UNWINDOWED_568 ,
										MUX_10_1_IN_9 => UNWINDOWED_57 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_540
									);
MUX_REORD_UNIT_541 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_541 ,
										MUX_10_1_IN_1 => UNWINDOWED_542 ,
										MUX_10_1_IN_2 => UNWINDOWED_539 ,
										MUX_10_1_IN_3 => UNWINDOWED_539 ,
										MUX_10_1_IN_4 => UNWINDOWED_539 ,
										MUX_10_1_IN_5 => UNWINDOWED_570 ,
										MUX_10_1_IN_6 => UNWINDOWED_570 ,
										MUX_10_1_IN_7 => UNWINDOWED_570 ,
										MUX_10_1_IN_8 => UNWINDOWED_570 ,
										MUX_10_1_IN_9 => UNWINDOWED_59 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_541
									);
MUX_REORD_UNIT_542 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_542 ,
										MUX_10_1_IN_1 => UNWINDOWED_541 ,
										MUX_10_1_IN_2 => UNWINDOWED_541 ,
										MUX_10_1_IN_3 => UNWINDOWED_541 ,
										MUX_10_1_IN_4 => UNWINDOWED_541 ,
										MUX_10_1_IN_5 => UNWINDOWED_572 ,
										MUX_10_1_IN_6 => UNWINDOWED_572 ,
										MUX_10_1_IN_7 => UNWINDOWED_572 ,
										MUX_10_1_IN_8 => UNWINDOWED_572 ,
										MUX_10_1_IN_9 => UNWINDOWED_61 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_542
									);
MUX_REORD_UNIT_543 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_543 ,
										MUX_10_1_IN_1 => UNWINDOWED_543 ,
										MUX_10_1_IN_2 => UNWINDOWED_543 ,
										MUX_10_1_IN_3 => UNWINDOWED_543 ,
										MUX_10_1_IN_4 => UNWINDOWED_543 ,
										MUX_10_1_IN_5 => UNWINDOWED_574 ,
										MUX_10_1_IN_6 => UNWINDOWED_574 ,
										MUX_10_1_IN_7 => UNWINDOWED_574 ,
										MUX_10_1_IN_8 => UNWINDOWED_574 ,
										MUX_10_1_IN_9 => UNWINDOWED_63 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_543
									);
MUX_REORD_UNIT_544 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_544 ,
										MUX_10_1_IN_1 => UNWINDOWED_544 ,
										MUX_10_1_IN_2 => UNWINDOWED_544 ,
										MUX_10_1_IN_3 => UNWINDOWED_544 ,
										MUX_10_1_IN_4 => UNWINDOWED_544 ,
										MUX_10_1_IN_5 => UNWINDOWED_513 ,
										MUX_10_1_IN_6 => UNWINDOWED_576 ,
										MUX_10_1_IN_7 => UNWINDOWED_576 ,
										MUX_10_1_IN_8 => UNWINDOWED_576 ,
										MUX_10_1_IN_9 => UNWINDOWED_65 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_544
									);
MUX_REORD_UNIT_545 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_545 ,
										MUX_10_1_IN_1 => UNWINDOWED_546 ,
										MUX_10_1_IN_2 => UNWINDOWED_546 ,
										MUX_10_1_IN_3 => UNWINDOWED_546 ,
										MUX_10_1_IN_4 => UNWINDOWED_546 ,
										MUX_10_1_IN_5 => UNWINDOWED_515 ,
										MUX_10_1_IN_6 => UNWINDOWED_578 ,
										MUX_10_1_IN_7 => UNWINDOWED_578 ,
										MUX_10_1_IN_8 => UNWINDOWED_578 ,
										MUX_10_1_IN_9 => UNWINDOWED_67 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_545
									);
MUX_REORD_UNIT_546 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_546 ,
										MUX_10_1_IN_1 => UNWINDOWED_545 ,
										MUX_10_1_IN_2 => UNWINDOWED_548 ,
										MUX_10_1_IN_3 => UNWINDOWED_548 ,
										MUX_10_1_IN_4 => UNWINDOWED_548 ,
										MUX_10_1_IN_5 => UNWINDOWED_517 ,
										MUX_10_1_IN_6 => UNWINDOWED_580 ,
										MUX_10_1_IN_7 => UNWINDOWED_580 ,
										MUX_10_1_IN_8 => UNWINDOWED_580 ,
										MUX_10_1_IN_9 => UNWINDOWED_69 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_546
									);
MUX_REORD_UNIT_547 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_547 ,
										MUX_10_1_IN_1 => UNWINDOWED_547 ,
										MUX_10_1_IN_2 => UNWINDOWED_550 ,
										MUX_10_1_IN_3 => UNWINDOWED_550 ,
										MUX_10_1_IN_4 => UNWINDOWED_550 ,
										MUX_10_1_IN_5 => UNWINDOWED_519 ,
										MUX_10_1_IN_6 => UNWINDOWED_582 ,
										MUX_10_1_IN_7 => UNWINDOWED_582 ,
										MUX_10_1_IN_8 => UNWINDOWED_582 ,
										MUX_10_1_IN_9 => UNWINDOWED_71 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_547
									);
MUX_REORD_UNIT_548 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_548 ,
										MUX_10_1_IN_1 => UNWINDOWED_548 ,
										MUX_10_1_IN_2 => UNWINDOWED_545 ,
										MUX_10_1_IN_3 => UNWINDOWED_552 ,
										MUX_10_1_IN_4 => UNWINDOWED_552 ,
										MUX_10_1_IN_5 => UNWINDOWED_521 ,
										MUX_10_1_IN_6 => UNWINDOWED_584 ,
										MUX_10_1_IN_7 => UNWINDOWED_584 ,
										MUX_10_1_IN_8 => UNWINDOWED_584 ,
										MUX_10_1_IN_9 => UNWINDOWED_73 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_548
									);
MUX_REORD_UNIT_549 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_549 ,
										MUX_10_1_IN_1 => UNWINDOWED_550 ,
										MUX_10_1_IN_2 => UNWINDOWED_547 ,
										MUX_10_1_IN_3 => UNWINDOWED_554 ,
										MUX_10_1_IN_4 => UNWINDOWED_554 ,
										MUX_10_1_IN_5 => UNWINDOWED_523 ,
										MUX_10_1_IN_6 => UNWINDOWED_586 ,
										MUX_10_1_IN_7 => UNWINDOWED_586 ,
										MUX_10_1_IN_8 => UNWINDOWED_586 ,
										MUX_10_1_IN_9 => UNWINDOWED_75 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_549
									);
MUX_REORD_UNIT_550 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_550 ,
										MUX_10_1_IN_1 => UNWINDOWED_549 ,
										MUX_10_1_IN_2 => UNWINDOWED_549 ,
										MUX_10_1_IN_3 => UNWINDOWED_556 ,
										MUX_10_1_IN_4 => UNWINDOWED_556 ,
										MUX_10_1_IN_5 => UNWINDOWED_525 ,
										MUX_10_1_IN_6 => UNWINDOWED_588 ,
										MUX_10_1_IN_7 => UNWINDOWED_588 ,
										MUX_10_1_IN_8 => UNWINDOWED_588 ,
										MUX_10_1_IN_9 => UNWINDOWED_77 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_550
									);
MUX_REORD_UNIT_551 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_551 ,
										MUX_10_1_IN_1 => UNWINDOWED_551 ,
										MUX_10_1_IN_2 => UNWINDOWED_551 ,
										MUX_10_1_IN_3 => UNWINDOWED_558 ,
										MUX_10_1_IN_4 => UNWINDOWED_558 ,
										MUX_10_1_IN_5 => UNWINDOWED_527 ,
										MUX_10_1_IN_6 => UNWINDOWED_590 ,
										MUX_10_1_IN_7 => UNWINDOWED_590 ,
										MUX_10_1_IN_8 => UNWINDOWED_590 ,
										MUX_10_1_IN_9 => UNWINDOWED_79 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_551
									);
MUX_REORD_UNIT_552 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_552 ,
										MUX_10_1_IN_1 => UNWINDOWED_552 ,
										MUX_10_1_IN_2 => UNWINDOWED_552 ,
										MUX_10_1_IN_3 => UNWINDOWED_545 ,
										MUX_10_1_IN_4 => UNWINDOWED_560 ,
										MUX_10_1_IN_5 => UNWINDOWED_529 ,
										MUX_10_1_IN_6 => UNWINDOWED_592 ,
										MUX_10_1_IN_7 => UNWINDOWED_592 ,
										MUX_10_1_IN_8 => UNWINDOWED_592 ,
										MUX_10_1_IN_9 => UNWINDOWED_81 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_552
									);
MUX_REORD_UNIT_553 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_553 ,
										MUX_10_1_IN_1 => UNWINDOWED_554 ,
										MUX_10_1_IN_2 => UNWINDOWED_554 ,
										MUX_10_1_IN_3 => UNWINDOWED_547 ,
										MUX_10_1_IN_4 => UNWINDOWED_562 ,
										MUX_10_1_IN_5 => UNWINDOWED_531 ,
										MUX_10_1_IN_6 => UNWINDOWED_594 ,
										MUX_10_1_IN_7 => UNWINDOWED_594 ,
										MUX_10_1_IN_8 => UNWINDOWED_594 ,
										MUX_10_1_IN_9 => UNWINDOWED_83 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_553
									);
MUX_REORD_UNIT_554 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_554 ,
										MUX_10_1_IN_1 => UNWINDOWED_553 ,
										MUX_10_1_IN_2 => UNWINDOWED_556 ,
										MUX_10_1_IN_3 => UNWINDOWED_549 ,
										MUX_10_1_IN_4 => UNWINDOWED_564 ,
										MUX_10_1_IN_5 => UNWINDOWED_533 ,
										MUX_10_1_IN_6 => UNWINDOWED_596 ,
										MUX_10_1_IN_7 => UNWINDOWED_596 ,
										MUX_10_1_IN_8 => UNWINDOWED_596 ,
										MUX_10_1_IN_9 => UNWINDOWED_85 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_554
									);
MUX_REORD_UNIT_555 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_555 ,
										MUX_10_1_IN_1 => UNWINDOWED_555 ,
										MUX_10_1_IN_2 => UNWINDOWED_558 ,
										MUX_10_1_IN_3 => UNWINDOWED_551 ,
										MUX_10_1_IN_4 => UNWINDOWED_566 ,
										MUX_10_1_IN_5 => UNWINDOWED_535 ,
										MUX_10_1_IN_6 => UNWINDOWED_598 ,
										MUX_10_1_IN_7 => UNWINDOWED_598 ,
										MUX_10_1_IN_8 => UNWINDOWED_598 ,
										MUX_10_1_IN_9 => UNWINDOWED_87 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_555
									);
MUX_REORD_UNIT_556 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_556 ,
										MUX_10_1_IN_1 => UNWINDOWED_556 ,
										MUX_10_1_IN_2 => UNWINDOWED_553 ,
										MUX_10_1_IN_3 => UNWINDOWED_553 ,
										MUX_10_1_IN_4 => UNWINDOWED_568 ,
										MUX_10_1_IN_5 => UNWINDOWED_537 ,
										MUX_10_1_IN_6 => UNWINDOWED_600 ,
										MUX_10_1_IN_7 => UNWINDOWED_600 ,
										MUX_10_1_IN_8 => UNWINDOWED_600 ,
										MUX_10_1_IN_9 => UNWINDOWED_89 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_556
									);
MUX_REORD_UNIT_557 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_557 ,
										MUX_10_1_IN_1 => UNWINDOWED_558 ,
										MUX_10_1_IN_2 => UNWINDOWED_555 ,
										MUX_10_1_IN_3 => UNWINDOWED_555 ,
										MUX_10_1_IN_4 => UNWINDOWED_570 ,
										MUX_10_1_IN_5 => UNWINDOWED_539 ,
										MUX_10_1_IN_6 => UNWINDOWED_602 ,
										MUX_10_1_IN_7 => UNWINDOWED_602 ,
										MUX_10_1_IN_8 => UNWINDOWED_602 ,
										MUX_10_1_IN_9 => UNWINDOWED_91 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_557
									);
MUX_REORD_UNIT_558 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_558 ,
										MUX_10_1_IN_1 => UNWINDOWED_557 ,
										MUX_10_1_IN_2 => UNWINDOWED_557 ,
										MUX_10_1_IN_3 => UNWINDOWED_557 ,
										MUX_10_1_IN_4 => UNWINDOWED_572 ,
										MUX_10_1_IN_5 => UNWINDOWED_541 ,
										MUX_10_1_IN_6 => UNWINDOWED_604 ,
										MUX_10_1_IN_7 => UNWINDOWED_604 ,
										MUX_10_1_IN_8 => UNWINDOWED_604 ,
										MUX_10_1_IN_9 => UNWINDOWED_93 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_558
									);
MUX_REORD_UNIT_559 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_559 ,
										MUX_10_1_IN_1 => UNWINDOWED_559 ,
										MUX_10_1_IN_2 => UNWINDOWED_559 ,
										MUX_10_1_IN_3 => UNWINDOWED_559 ,
										MUX_10_1_IN_4 => UNWINDOWED_574 ,
										MUX_10_1_IN_5 => UNWINDOWED_543 ,
										MUX_10_1_IN_6 => UNWINDOWED_606 ,
										MUX_10_1_IN_7 => UNWINDOWED_606 ,
										MUX_10_1_IN_8 => UNWINDOWED_606 ,
										MUX_10_1_IN_9 => UNWINDOWED_95 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_559
									);
MUX_REORD_UNIT_560 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_560 ,
										MUX_10_1_IN_1 => UNWINDOWED_560 ,
										MUX_10_1_IN_2 => UNWINDOWED_560 ,
										MUX_10_1_IN_3 => UNWINDOWED_560 ,
										MUX_10_1_IN_4 => UNWINDOWED_545 ,
										MUX_10_1_IN_5 => UNWINDOWED_545 ,
										MUX_10_1_IN_6 => UNWINDOWED_608 ,
										MUX_10_1_IN_7 => UNWINDOWED_608 ,
										MUX_10_1_IN_8 => UNWINDOWED_608 ,
										MUX_10_1_IN_9 => UNWINDOWED_97 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_560
									);
MUX_REORD_UNIT_561 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_561 ,
										MUX_10_1_IN_1 => UNWINDOWED_562 ,
										MUX_10_1_IN_2 => UNWINDOWED_562 ,
										MUX_10_1_IN_3 => UNWINDOWED_562 ,
										MUX_10_1_IN_4 => UNWINDOWED_547 ,
										MUX_10_1_IN_5 => UNWINDOWED_547 ,
										MUX_10_1_IN_6 => UNWINDOWED_610 ,
										MUX_10_1_IN_7 => UNWINDOWED_610 ,
										MUX_10_1_IN_8 => UNWINDOWED_610 ,
										MUX_10_1_IN_9 => UNWINDOWED_99 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_561
									);
MUX_REORD_UNIT_562 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_562 ,
										MUX_10_1_IN_1 => UNWINDOWED_561 ,
										MUX_10_1_IN_2 => UNWINDOWED_564 ,
										MUX_10_1_IN_3 => UNWINDOWED_564 ,
										MUX_10_1_IN_4 => UNWINDOWED_549 ,
										MUX_10_1_IN_5 => UNWINDOWED_549 ,
										MUX_10_1_IN_6 => UNWINDOWED_612 ,
										MUX_10_1_IN_7 => UNWINDOWED_612 ,
										MUX_10_1_IN_8 => UNWINDOWED_612 ,
										MUX_10_1_IN_9 => UNWINDOWED_101 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_562
									);
MUX_REORD_UNIT_563 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_563 ,
										MUX_10_1_IN_1 => UNWINDOWED_563 ,
										MUX_10_1_IN_2 => UNWINDOWED_566 ,
										MUX_10_1_IN_3 => UNWINDOWED_566 ,
										MUX_10_1_IN_4 => UNWINDOWED_551 ,
										MUX_10_1_IN_5 => UNWINDOWED_551 ,
										MUX_10_1_IN_6 => UNWINDOWED_614 ,
										MUX_10_1_IN_7 => UNWINDOWED_614 ,
										MUX_10_1_IN_8 => UNWINDOWED_614 ,
										MUX_10_1_IN_9 => UNWINDOWED_103 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_563
									);
MUX_REORD_UNIT_564 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_564 ,
										MUX_10_1_IN_1 => UNWINDOWED_564 ,
										MUX_10_1_IN_2 => UNWINDOWED_561 ,
										MUX_10_1_IN_3 => UNWINDOWED_568 ,
										MUX_10_1_IN_4 => UNWINDOWED_553 ,
										MUX_10_1_IN_5 => UNWINDOWED_553 ,
										MUX_10_1_IN_6 => UNWINDOWED_616 ,
										MUX_10_1_IN_7 => UNWINDOWED_616 ,
										MUX_10_1_IN_8 => UNWINDOWED_616 ,
										MUX_10_1_IN_9 => UNWINDOWED_105 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_564
									);
MUX_REORD_UNIT_565 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_565 ,
										MUX_10_1_IN_1 => UNWINDOWED_566 ,
										MUX_10_1_IN_2 => UNWINDOWED_563 ,
										MUX_10_1_IN_3 => UNWINDOWED_570 ,
										MUX_10_1_IN_4 => UNWINDOWED_555 ,
										MUX_10_1_IN_5 => UNWINDOWED_555 ,
										MUX_10_1_IN_6 => UNWINDOWED_618 ,
										MUX_10_1_IN_7 => UNWINDOWED_618 ,
										MUX_10_1_IN_8 => UNWINDOWED_618 ,
										MUX_10_1_IN_9 => UNWINDOWED_107 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_565
									);
MUX_REORD_UNIT_566 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_566 ,
										MUX_10_1_IN_1 => UNWINDOWED_565 ,
										MUX_10_1_IN_2 => UNWINDOWED_565 ,
										MUX_10_1_IN_3 => UNWINDOWED_572 ,
										MUX_10_1_IN_4 => UNWINDOWED_557 ,
										MUX_10_1_IN_5 => UNWINDOWED_557 ,
										MUX_10_1_IN_6 => UNWINDOWED_620 ,
										MUX_10_1_IN_7 => UNWINDOWED_620 ,
										MUX_10_1_IN_8 => UNWINDOWED_620 ,
										MUX_10_1_IN_9 => UNWINDOWED_109 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_566
									);
MUX_REORD_UNIT_567 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_567 ,
										MUX_10_1_IN_1 => UNWINDOWED_567 ,
										MUX_10_1_IN_2 => UNWINDOWED_567 ,
										MUX_10_1_IN_3 => UNWINDOWED_574 ,
										MUX_10_1_IN_4 => UNWINDOWED_559 ,
										MUX_10_1_IN_5 => UNWINDOWED_559 ,
										MUX_10_1_IN_6 => UNWINDOWED_622 ,
										MUX_10_1_IN_7 => UNWINDOWED_622 ,
										MUX_10_1_IN_8 => UNWINDOWED_622 ,
										MUX_10_1_IN_9 => UNWINDOWED_111 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_567
									);
MUX_REORD_UNIT_568 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_568 ,
										MUX_10_1_IN_1 => UNWINDOWED_568 ,
										MUX_10_1_IN_2 => UNWINDOWED_568 ,
										MUX_10_1_IN_3 => UNWINDOWED_561 ,
										MUX_10_1_IN_4 => UNWINDOWED_561 ,
										MUX_10_1_IN_5 => UNWINDOWED_561 ,
										MUX_10_1_IN_6 => UNWINDOWED_624 ,
										MUX_10_1_IN_7 => UNWINDOWED_624 ,
										MUX_10_1_IN_8 => UNWINDOWED_624 ,
										MUX_10_1_IN_9 => UNWINDOWED_113 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_568
									);
MUX_REORD_UNIT_569 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_569 ,
										MUX_10_1_IN_1 => UNWINDOWED_570 ,
										MUX_10_1_IN_2 => UNWINDOWED_570 ,
										MUX_10_1_IN_3 => UNWINDOWED_563 ,
										MUX_10_1_IN_4 => UNWINDOWED_563 ,
										MUX_10_1_IN_5 => UNWINDOWED_563 ,
										MUX_10_1_IN_6 => UNWINDOWED_626 ,
										MUX_10_1_IN_7 => UNWINDOWED_626 ,
										MUX_10_1_IN_8 => UNWINDOWED_626 ,
										MUX_10_1_IN_9 => UNWINDOWED_115 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_569
									);
MUX_REORD_UNIT_570 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_570 ,
										MUX_10_1_IN_1 => UNWINDOWED_569 ,
										MUX_10_1_IN_2 => UNWINDOWED_572 ,
										MUX_10_1_IN_3 => UNWINDOWED_565 ,
										MUX_10_1_IN_4 => UNWINDOWED_565 ,
										MUX_10_1_IN_5 => UNWINDOWED_565 ,
										MUX_10_1_IN_6 => UNWINDOWED_628 ,
										MUX_10_1_IN_7 => UNWINDOWED_628 ,
										MUX_10_1_IN_8 => UNWINDOWED_628 ,
										MUX_10_1_IN_9 => UNWINDOWED_117 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_570
									);
MUX_REORD_UNIT_571 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_571 ,
										MUX_10_1_IN_1 => UNWINDOWED_571 ,
										MUX_10_1_IN_2 => UNWINDOWED_574 ,
										MUX_10_1_IN_3 => UNWINDOWED_567 ,
										MUX_10_1_IN_4 => UNWINDOWED_567 ,
										MUX_10_1_IN_5 => UNWINDOWED_567 ,
										MUX_10_1_IN_6 => UNWINDOWED_630 ,
										MUX_10_1_IN_7 => UNWINDOWED_630 ,
										MUX_10_1_IN_8 => UNWINDOWED_630 ,
										MUX_10_1_IN_9 => UNWINDOWED_119 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_571
									);
MUX_REORD_UNIT_572 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_572 ,
										MUX_10_1_IN_1 => UNWINDOWED_572 ,
										MUX_10_1_IN_2 => UNWINDOWED_569 ,
										MUX_10_1_IN_3 => UNWINDOWED_569 ,
										MUX_10_1_IN_4 => UNWINDOWED_569 ,
										MUX_10_1_IN_5 => UNWINDOWED_569 ,
										MUX_10_1_IN_6 => UNWINDOWED_632 ,
										MUX_10_1_IN_7 => UNWINDOWED_632 ,
										MUX_10_1_IN_8 => UNWINDOWED_632 ,
										MUX_10_1_IN_9 => UNWINDOWED_121 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_572
									);
MUX_REORD_UNIT_573 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_573 ,
										MUX_10_1_IN_1 => UNWINDOWED_574 ,
										MUX_10_1_IN_2 => UNWINDOWED_571 ,
										MUX_10_1_IN_3 => UNWINDOWED_571 ,
										MUX_10_1_IN_4 => UNWINDOWED_571 ,
										MUX_10_1_IN_5 => UNWINDOWED_571 ,
										MUX_10_1_IN_6 => UNWINDOWED_634 ,
										MUX_10_1_IN_7 => UNWINDOWED_634 ,
										MUX_10_1_IN_8 => UNWINDOWED_634 ,
										MUX_10_1_IN_9 => UNWINDOWED_123 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_573
									);
MUX_REORD_UNIT_574 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_574 ,
										MUX_10_1_IN_1 => UNWINDOWED_573 ,
										MUX_10_1_IN_2 => UNWINDOWED_573 ,
										MUX_10_1_IN_3 => UNWINDOWED_573 ,
										MUX_10_1_IN_4 => UNWINDOWED_573 ,
										MUX_10_1_IN_5 => UNWINDOWED_573 ,
										MUX_10_1_IN_6 => UNWINDOWED_636 ,
										MUX_10_1_IN_7 => UNWINDOWED_636 ,
										MUX_10_1_IN_8 => UNWINDOWED_636 ,
										MUX_10_1_IN_9 => UNWINDOWED_125 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_574
									);
MUX_REORD_UNIT_575 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_575 ,
										MUX_10_1_IN_1 => UNWINDOWED_575 ,
										MUX_10_1_IN_2 => UNWINDOWED_575 ,
										MUX_10_1_IN_3 => UNWINDOWED_575 ,
										MUX_10_1_IN_4 => UNWINDOWED_575 ,
										MUX_10_1_IN_5 => UNWINDOWED_575 ,
										MUX_10_1_IN_6 => UNWINDOWED_638 ,
										MUX_10_1_IN_7 => UNWINDOWED_638 ,
										MUX_10_1_IN_8 => UNWINDOWED_638 ,
										MUX_10_1_IN_9 => UNWINDOWED_127 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_575
									);
MUX_REORD_UNIT_576 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_576 ,
										MUX_10_1_IN_1 => UNWINDOWED_576 ,
										MUX_10_1_IN_2 => UNWINDOWED_576 ,
										MUX_10_1_IN_3 => UNWINDOWED_576 ,
										MUX_10_1_IN_4 => UNWINDOWED_576 ,
										MUX_10_1_IN_5 => UNWINDOWED_576 ,
										MUX_10_1_IN_6 => UNWINDOWED_513 ,
										MUX_10_1_IN_7 => UNWINDOWED_640 ,
										MUX_10_1_IN_8 => UNWINDOWED_640 ,
										MUX_10_1_IN_9 => UNWINDOWED_129 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_576
									);
MUX_REORD_UNIT_577 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_577 ,
										MUX_10_1_IN_1 => UNWINDOWED_578 ,
										MUX_10_1_IN_2 => UNWINDOWED_578 ,
										MUX_10_1_IN_3 => UNWINDOWED_578 ,
										MUX_10_1_IN_4 => UNWINDOWED_578 ,
										MUX_10_1_IN_5 => UNWINDOWED_578 ,
										MUX_10_1_IN_6 => UNWINDOWED_515 ,
										MUX_10_1_IN_7 => UNWINDOWED_642 ,
										MUX_10_1_IN_8 => UNWINDOWED_642 ,
										MUX_10_1_IN_9 => UNWINDOWED_131 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_577
									);
MUX_REORD_UNIT_578 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_578 ,
										MUX_10_1_IN_1 => UNWINDOWED_577 ,
										MUX_10_1_IN_2 => UNWINDOWED_580 ,
										MUX_10_1_IN_3 => UNWINDOWED_580 ,
										MUX_10_1_IN_4 => UNWINDOWED_580 ,
										MUX_10_1_IN_5 => UNWINDOWED_580 ,
										MUX_10_1_IN_6 => UNWINDOWED_517 ,
										MUX_10_1_IN_7 => UNWINDOWED_644 ,
										MUX_10_1_IN_8 => UNWINDOWED_644 ,
										MUX_10_1_IN_9 => UNWINDOWED_133 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_578
									);
MUX_REORD_UNIT_579 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_579 ,
										MUX_10_1_IN_1 => UNWINDOWED_579 ,
										MUX_10_1_IN_2 => UNWINDOWED_582 ,
										MUX_10_1_IN_3 => UNWINDOWED_582 ,
										MUX_10_1_IN_4 => UNWINDOWED_582 ,
										MUX_10_1_IN_5 => UNWINDOWED_582 ,
										MUX_10_1_IN_6 => UNWINDOWED_519 ,
										MUX_10_1_IN_7 => UNWINDOWED_646 ,
										MUX_10_1_IN_8 => UNWINDOWED_646 ,
										MUX_10_1_IN_9 => UNWINDOWED_135 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_579
									);
MUX_REORD_UNIT_580 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_580 ,
										MUX_10_1_IN_1 => UNWINDOWED_580 ,
										MUX_10_1_IN_2 => UNWINDOWED_577 ,
										MUX_10_1_IN_3 => UNWINDOWED_584 ,
										MUX_10_1_IN_4 => UNWINDOWED_584 ,
										MUX_10_1_IN_5 => UNWINDOWED_584 ,
										MUX_10_1_IN_6 => UNWINDOWED_521 ,
										MUX_10_1_IN_7 => UNWINDOWED_648 ,
										MUX_10_1_IN_8 => UNWINDOWED_648 ,
										MUX_10_1_IN_9 => UNWINDOWED_137 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_580
									);
MUX_REORD_UNIT_581 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_581 ,
										MUX_10_1_IN_1 => UNWINDOWED_582 ,
										MUX_10_1_IN_2 => UNWINDOWED_579 ,
										MUX_10_1_IN_3 => UNWINDOWED_586 ,
										MUX_10_1_IN_4 => UNWINDOWED_586 ,
										MUX_10_1_IN_5 => UNWINDOWED_586 ,
										MUX_10_1_IN_6 => UNWINDOWED_523 ,
										MUX_10_1_IN_7 => UNWINDOWED_650 ,
										MUX_10_1_IN_8 => UNWINDOWED_650 ,
										MUX_10_1_IN_9 => UNWINDOWED_139 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_581
									);
MUX_REORD_UNIT_582 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_582 ,
										MUX_10_1_IN_1 => UNWINDOWED_581 ,
										MUX_10_1_IN_2 => UNWINDOWED_581 ,
										MUX_10_1_IN_3 => UNWINDOWED_588 ,
										MUX_10_1_IN_4 => UNWINDOWED_588 ,
										MUX_10_1_IN_5 => UNWINDOWED_588 ,
										MUX_10_1_IN_6 => UNWINDOWED_525 ,
										MUX_10_1_IN_7 => UNWINDOWED_652 ,
										MUX_10_1_IN_8 => UNWINDOWED_652 ,
										MUX_10_1_IN_9 => UNWINDOWED_141 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_582
									);
MUX_REORD_UNIT_583 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_583 ,
										MUX_10_1_IN_1 => UNWINDOWED_583 ,
										MUX_10_1_IN_2 => UNWINDOWED_583 ,
										MUX_10_1_IN_3 => UNWINDOWED_590 ,
										MUX_10_1_IN_4 => UNWINDOWED_590 ,
										MUX_10_1_IN_5 => UNWINDOWED_590 ,
										MUX_10_1_IN_6 => UNWINDOWED_527 ,
										MUX_10_1_IN_7 => UNWINDOWED_654 ,
										MUX_10_1_IN_8 => UNWINDOWED_654 ,
										MUX_10_1_IN_9 => UNWINDOWED_143 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_583
									);
MUX_REORD_UNIT_584 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_584 ,
										MUX_10_1_IN_1 => UNWINDOWED_584 ,
										MUX_10_1_IN_2 => UNWINDOWED_584 ,
										MUX_10_1_IN_3 => UNWINDOWED_577 ,
										MUX_10_1_IN_4 => UNWINDOWED_592 ,
										MUX_10_1_IN_5 => UNWINDOWED_592 ,
										MUX_10_1_IN_6 => UNWINDOWED_529 ,
										MUX_10_1_IN_7 => UNWINDOWED_656 ,
										MUX_10_1_IN_8 => UNWINDOWED_656 ,
										MUX_10_1_IN_9 => UNWINDOWED_145 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_584
									);
MUX_REORD_UNIT_585 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_585 ,
										MUX_10_1_IN_1 => UNWINDOWED_586 ,
										MUX_10_1_IN_2 => UNWINDOWED_586 ,
										MUX_10_1_IN_3 => UNWINDOWED_579 ,
										MUX_10_1_IN_4 => UNWINDOWED_594 ,
										MUX_10_1_IN_5 => UNWINDOWED_594 ,
										MUX_10_1_IN_6 => UNWINDOWED_531 ,
										MUX_10_1_IN_7 => UNWINDOWED_658 ,
										MUX_10_1_IN_8 => UNWINDOWED_658 ,
										MUX_10_1_IN_9 => UNWINDOWED_147 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_585
									);
MUX_REORD_UNIT_586 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_586 ,
										MUX_10_1_IN_1 => UNWINDOWED_585 ,
										MUX_10_1_IN_2 => UNWINDOWED_588 ,
										MUX_10_1_IN_3 => UNWINDOWED_581 ,
										MUX_10_1_IN_4 => UNWINDOWED_596 ,
										MUX_10_1_IN_5 => UNWINDOWED_596 ,
										MUX_10_1_IN_6 => UNWINDOWED_533 ,
										MUX_10_1_IN_7 => UNWINDOWED_660 ,
										MUX_10_1_IN_8 => UNWINDOWED_660 ,
										MUX_10_1_IN_9 => UNWINDOWED_149 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_586
									);
MUX_REORD_UNIT_587 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_587 ,
										MUX_10_1_IN_1 => UNWINDOWED_587 ,
										MUX_10_1_IN_2 => UNWINDOWED_590 ,
										MUX_10_1_IN_3 => UNWINDOWED_583 ,
										MUX_10_1_IN_4 => UNWINDOWED_598 ,
										MUX_10_1_IN_5 => UNWINDOWED_598 ,
										MUX_10_1_IN_6 => UNWINDOWED_535 ,
										MUX_10_1_IN_7 => UNWINDOWED_662 ,
										MUX_10_1_IN_8 => UNWINDOWED_662 ,
										MUX_10_1_IN_9 => UNWINDOWED_151 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_587
									);
MUX_REORD_UNIT_588 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_588 ,
										MUX_10_1_IN_1 => UNWINDOWED_588 ,
										MUX_10_1_IN_2 => UNWINDOWED_585 ,
										MUX_10_1_IN_3 => UNWINDOWED_585 ,
										MUX_10_1_IN_4 => UNWINDOWED_600 ,
										MUX_10_1_IN_5 => UNWINDOWED_600 ,
										MUX_10_1_IN_6 => UNWINDOWED_537 ,
										MUX_10_1_IN_7 => UNWINDOWED_664 ,
										MUX_10_1_IN_8 => UNWINDOWED_664 ,
										MUX_10_1_IN_9 => UNWINDOWED_153 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_588
									);
MUX_REORD_UNIT_589 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_589 ,
										MUX_10_1_IN_1 => UNWINDOWED_590 ,
										MUX_10_1_IN_2 => UNWINDOWED_587 ,
										MUX_10_1_IN_3 => UNWINDOWED_587 ,
										MUX_10_1_IN_4 => UNWINDOWED_602 ,
										MUX_10_1_IN_5 => UNWINDOWED_602 ,
										MUX_10_1_IN_6 => UNWINDOWED_539 ,
										MUX_10_1_IN_7 => UNWINDOWED_666 ,
										MUX_10_1_IN_8 => UNWINDOWED_666 ,
										MUX_10_1_IN_9 => UNWINDOWED_155 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_589
									);
MUX_REORD_UNIT_590 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_590 ,
										MUX_10_1_IN_1 => UNWINDOWED_589 ,
										MUX_10_1_IN_2 => UNWINDOWED_589 ,
										MUX_10_1_IN_3 => UNWINDOWED_589 ,
										MUX_10_1_IN_4 => UNWINDOWED_604 ,
										MUX_10_1_IN_5 => UNWINDOWED_604 ,
										MUX_10_1_IN_6 => UNWINDOWED_541 ,
										MUX_10_1_IN_7 => UNWINDOWED_668 ,
										MUX_10_1_IN_8 => UNWINDOWED_668 ,
										MUX_10_1_IN_9 => UNWINDOWED_157 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_590
									);
MUX_REORD_UNIT_591 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_591 ,
										MUX_10_1_IN_1 => UNWINDOWED_591 ,
										MUX_10_1_IN_2 => UNWINDOWED_591 ,
										MUX_10_1_IN_3 => UNWINDOWED_591 ,
										MUX_10_1_IN_4 => UNWINDOWED_606 ,
										MUX_10_1_IN_5 => UNWINDOWED_606 ,
										MUX_10_1_IN_6 => UNWINDOWED_543 ,
										MUX_10_1_IN_7 => UNWINDOWED_670 ,
										MUX_10_1_IN_8 => UNWINDOWED_670 ,
										MUX_10_1_IN_9 => UNWINDOWED_159 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_591
									);
MUX_REORD_UNIT_592 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_592 ,
										MUX_10_1_IN_1 => UNWINDOWED_592 ,
										MUX_10_1_IN_2 => UNWINDOWED_592 ,
										MUX_10_1_IN_3 => UNWINDOWED_592 ,
										MUX_10_1_IN_4 => UNWINDOWED_577 ,
										MUX_10_1_IN_5 => UNWINDOWED_608 ,
										MUX_10_1_IN_6 => UNWINDOWED_545 ,
										MUX_10_1_IN_7 => UNWINDOWED_672 ,
										MUX_10_1_IN_8 => UNWINDOWED_672 ,
										MUX_10_1_IN_9 => UNWINDOWED_161 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_592
									);
MUX_REORD_UNIT_593 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_593 ,
										MUX_10_1_IN_1 => UNWINDOWED_594 ,
										MUX_10_1_IN_2 => UNWINDOWED_594 ,
										MUX_10_1_IN_3 => UNWINDOWED_594 ,
										MUX_10_1_IN_4 => UNWINDOWED_579 ,
										MUX_10_1_IN_5 => UNWINDOWED_610 ,
										MUX_10_1_IN_6 => UNWINDOWED_547 ,
										MUX_10_1_IN_7 => UNWINDOWED_674 ,
										MUX_10_1_IN_8 => UNWINDOWED_674 ,
										MUX_10_1_IN_9 => UNWINDOWED_163 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_593
									);
MUX_REORD_UNIT_594 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_594 ,
										MUX_10_1_IN_1 => UNWINDOWED_593 ,
										MUX_10_1_IN_2 => UNWINDOWED_596 ,
										MUX_10_1_IN_3 => UNWINDOWED_596 ,
										MUX_10_1_IN_4 => UNWINDOWED_581 ,
										MUX_10_1_IN_5 => UNWINDOWED_612 ,
										MUX_10_1_IN_6 => UNWINDOWED_549 ,
										MUX_10_1_IN_7 => UNWINDOWED_676 ,
										MUX_10_1_IN_8 => UNWINDOWED_676 ,
										MUX_10_1_IN_9 => UNWINDOWED_165 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_594
									);
MUX_REORD_UNIT_595 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_595 ,
										MUX_10_1_IN_1 => UNWINDOWED_595 ,
										MUX_10_1_IN_2 => UNWINDOWED_598 ,
										MUX_10_1_IN_3 => UNWINDOWED_598 ,
										MUX_10_1_IN_4 => UNWINDOWED_583 ,
										MUX_10_1_IN_5 => UNWINDOWED_614 ,
										MUX_10_1_IN_6 => UNWINDOWED_551 ,
										MUX_10_1_IN_7 => UNWINDOWED_678 ,
										MUX_10_1_IN_8 => UNWINDOWED_678 ,
										MUX_10_1_IN_9 => UNWINDOWED_167 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_595
									);
MUX_REORD_UNIT_596 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_596 ,
										MUX_10_1_IN_1 => UNWINDOWED_596 ,
										MUX_10_1_IN_2 => UNWINDOWED_593 ,
										MUX_10_1_IN_3 => UNWINDOWED_600 ,
										MUX_10_1_IN_4 => UNWINDOWED_585 ,
										MUX_10_1_IN_5 => UNWINDOWED_616 ,
										MUX_10_1_IN_6 => UNWINDOWED_553 ,
										MUX_10_1_IN_7 => UNWINDOWED_680 ,
										MUX_10_1_IN_8 => UNWINDOWED_680 ,
										MUX_10_1_IN_9 => UNWINDOWED_169 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_596
									);
MUX_REORD_UNIT_597 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_597 ,
										MUX_10_1_IN_1 => UNWINDOWED_598 ,
										MUX_10_1_IN_2 => UNWINDOWED_595 ,
										MUX_10_1_IN_3 => UNWINDOWED_602 ,
										MUX_10_1_IN_4 => UNWINDOWED_587 ,
										MUX_10_1_IN_5 => UNWINDOWED_618 ,
										MUX_10_1_IN_6 => UNWINDOWED_555 ,
										MUX_10_1_IN_7 => UNWINDOWED_682 ,
										MUX_10_1_IN_8 => UNWINDOWED_682 ,
										MUX_10_1_IN_9 => UNWINDOWED_171 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_597
									);
MUX_REORD_UNIT_598 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_598 ,
										MUX_10_1_IN_1 => UNWINDOWED_597 ,
										MUX_10_1_IN_2 => UNWINDOWED_597 ,
										MUX_10_1_IN_3 => UNWINDOWED_604 ,
										MUX_10_1_IN_4 => UNWINDOWED_589 ,
										MUX_10_1_IN_5 => UNWINDOWED_620 ,
										MUX_10_1_IN_6 => UNWINDOWED_557 ,
										MUX_10_1_IN_7 => UNWINDOWED_684 ,
										MUX_10_1_IN_8 => UNWINDOWED_684 ,
										MUX_10_1_IN_9 => UNWINDOWED_173 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_598
									);
MUX_REORD_UNIT_599 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_599 ,
										MUX_10_1_IN_1 => UNWINDOWED_599 ,
										MUX_10_1_IN_2 => UNWINDOWED_599 ,
										MUX_10_1_IN_3 => UNWINDOWED_606 ,
										MUX_10_1_IN_4 => UNWINDOWED_591 ,
										MUX_10_1_IN_5 => UNWINDOWED_622 ,
										MUX_10_1_IN_6 => UNWINDOWED_559 ,
										MUX_10_1_IN_7 => UNWINDOWED_686 ,
										MUX_10_1_IN_8 => UNWINDOWED_686 ,
										MUX_10_1_IN_9 => UNWINDOWED_175 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_599
									);
MUX_REORD_UNIT_600 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_600 ,
										MUX_10_1_IN_1 => UNWINDOWED_600 ,
										MUX_10_1_IN_2 => UNWINDOWED_600 ,
										MUX_10_1_IN_3 => UNWINDOWED_593 ,
										MUX_10_1_IN_4 => UNWINDOWED_593 ,
										MUX_10_1_IN_5 => UNWINDOWED_624 ,
										MUX_10_1_IN_6 => UNWINDOWED_561 ,
										MUX_10_1_IN_7 => UNWINDOWED_688 ,
										MUX_10_1_IN_8 => UNWINDOWED_688 ,
										MUX_10_1_IN_9 => UNWINDOWED_177 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_600
									);
MUX_REORD_UNIT_601 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_601 ,
										MUX_10_1_IN_1 => UNWINDOWED_602 ,
										MUX_10_1_IN_2 => UNWINDOWED_602 ,
										MUX_10_1_IN_3 => UNWINDOWED_595 ,
										MUX_10_1_IN_4 => UNWINDOWED_595 ,
										MUX_10_1_IN_5 => UNWINDOWED_626 ,
										MUX_10_1_IN_6 => UNWINDOWED_563 ,
										MUX_10_1_IN_7 => UNWINDOWED_690 ,
										MUX_10_1_IN_8 => UNWINDOWED_690 ,
										MUX_10_1_IN_9 => UNWINDOWED_179 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_601
									);
MUX_REORD_UNIT_602 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_602 ,
										MUX_10_1_IN_1 => UNWINDOWED_601 ,
										MUX_10_1_IN_2 => UNWINDOWED_604 ,
										MUX_10_1_IN_3 => UNWINDOWED_597 ,
										MUX_10_1_IN_4 => UNWINDOWED_597 ,
										MUX_10_1_IN_5 => UNWINDOWED_628 ,
										MUX_10_1_IN_6 => UNWINDOWED_565 ,
										MUX_10_1_IN_7 => UNWINDOWED_692 ,
										MUX_10_1_IN_8 => UNWINDOWED_692 ,
										MUX_10_1_IN_9 => UNWINDOWED_181 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_602
									);
MUX_REORD_UNIT_603 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_603 ,
										MUX_10_1_IN_1 => UNWINDOWED_603 ,
										MUX_10_1_IN_2 => UNWINDOWED_606 ,
										MUX_10_1_IN_3 => UNWINDOWED_599 ,
										MUX_10_1_IN_4 => UNWINDOWED_599 ,
										MUX_10_1_IN_5 => UNWINDOWED_630 ,
										MUX_10_1_IN_6 => UNWINDOWED_567 ,
										MUX_10_1_IN_7 => UNWINDOWED_694 ,
										MUX_10_1_IN_8 => UNWINDOWED_694 ,
										MUX_10_1_IN_9 => UNWINDOWED_183 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_603
									);
MUX_REORD_UNIT_604 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_604 ,
										MUX_10_1_IN_1 => UNWINDOWED_604 ,
										MUX_10_1_IN_2 => UNWINDOWED_601 ,
										MUX_10_1_IN_3 => UNWINDOWED_601 ,
										MUX_10_1_IN_4 => UNWINDOWED_601 ,
										MUX_10_1_IN_5 => UNWINDOWED_632 ,
										MUX_10_1_IN_6 => UNWINDOWED_569 ,
										MUX_10_1_IN_7 => UNWINDOWED_696 ,
										MUX_10_1_IN_8 => UNWINDOWED_696 ,
										MUX_10_1_IN_9 => UNWINDOWED_185 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_604
									);
MUX_REORD_UNIT_605 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_605 ,
										MUX_10_1_IN_1 => UNWINDOWED_606 ,
										MUX_10_1_IN_2 => UNWINDOWED_603 ,
										MUX_10_1_IN_3 => UNWINDOWED_603 ,
										MUX_10_1_IN_4 => UNWINDOWED_603 ,
										MUX_10_1_IN_5 => UNWINDOWED_634 ,
										MUX_10_1_IN_6 => UNWINDOWED_571 ,
										MUX_10_1_IN_7 => UNWINDOWED_698 ,
										MUX_10_1_IN_8 => UNWINDOWED_698 ,
										MUX_10_1_IN_9 => UNWINDOWED_187 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_605
									);
MUX_REORD_UNIT_606 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_606 ,
										MUX_10_1_IN_1 => UNWINDOWED_605 ,
										MUX_10_1_IN_2 => UNWINDOWED_605 ,
										MUX_10_1_IN_3 => UNWINDOWED_605 ,
										MUX_10_1_IN_4 => UNWINDOWED_605 ,
										MUX_10_1_IN_5 => UNWINDOWED_636 ,
										MUX_10_1_IN_6 => UNWINDOWED_573 ,
										MUX_10_1_IN_7 => UNWINDOWED_700 ,
										MUX_10_1_IN_8 => UNWINDOWED_700 ,
										MUX_10_1_IN_9 => UNWINDOWED_189 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_606
									);
MUX_REORD_UNIT_607 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_607 ,
										MUX_10_1_IN_1 => UNWINDOWED_607 ,
										MUX_10_1_IN_2 => UNWINDOWED_607 ,
										MUX_10_1_IN_3 => UNWINDOWED_607 ,
										MUX_10_1_IN_4 => UNWINDOWED_607 ,
										MUX_10_1_IN_5 => UNWINDOWED_638 ,
										MUX_10_1_IN_6 => UNWINDOWED_575 ,
										MUX_10_1_IN_7 => UNWINDOWED_702 ,
										MUX_10_1_IN_8 => UNWINDOWED_702 ,
										MUX_10_1_IN_9 => UNWINDOWED_191 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_607
									);
MUX_REORD_UNIT_608 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_608 ,
										MUX_10_1_IN_1 => UNWINDOWED_608 ,
										MUX_10_1_IN_2 => UNWINDOWED_608 ,
										MUX_10_1_IN_3 => UNWINDOWED_608 ,
										MUX_10_1_IN_4 => UNWINDOWED_608 ,
										MUX_10_1_IN_5 => UNWINDOWED_577 ,
										MUX_10_1_IN_6 => UNWINDOWED_577 ,
										MUX_10_1_IN_7 => UNWINDOWED_704 ,
										MUX_10_1_IN_8 => UNWINDOWED_704 ,
										MUX_10_1_IN_9 => UNWINDOWED_193 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_608
									);
MUX_REORD_UNIT_609 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_609 ,
										MUX_10_1_IN_1 => UNWINDOWED_610 ,
										MUX_10_1_IN_2 => UNWINDOWED_610 ,
										MUX_10_1_IN_3 => UNWINDOWED_610 ,
										MUX_10_1_IN_4 => UNWINDOWED_610 ,
										MUX_10_1_IN_5 => UNWINDOWED_579 ,
										MUX_10_1_IN_6 => UNWINDOWED_579 ,
										MUX_10_1_IN_7 => UNWINDOWED_706 ,
										MUX_10_1_IN_8 => UNWINDOWED_706 ,
										MUX_10_1_IN_9 => UNWINDOWED_195 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_609
									);
MUX_REORD_UNIT_610 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_610 ,
										MUX_10_1_IN_1 => UNWINDOWED_609 ,
										MUX_10_1_IN_2 => UNWINDOWED_612 ,
										MUX_10_1_IN_3 => UNWINDOWED_612 ,
										MUX_10_1_IN_4 => UNWINDOWED_612 ,
										MUX_10_1_IN_5 => UNWINDOWED_581 ,
										MUX_10_1_IN_6 => UNWINDOWED_581 ,
										MUX_10_1_IN_7 => UNWINDOWED_708 ,
										MUX_10_1_IN_8 => UNWINDOWED_708 ,
										MUX_10_1_IN_9 => UNWINDOWED_197 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_610
									);
MUX_REORD_UNIT_611 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_611 ,
										MUX_10_1_IN_1 => UNWINDOWED_611 ,
										MUX_10_1_IN_2 => UNWINDOWED_614 ,
										MUX_10_1_IN_3 => UNWINDOWED_614 ,
										MUX_10_1_IN_4 => UNWINDOWED_614 ,
										MUX_10_1_IN_5 => UNWINDOWED_583 ,
										MUX_10_1_IN_6 => UNWINDOWED_583 ,
										MUX_10_1_IN_7 => UNWINDOWED_710 ,
										MUX_10_1_IN_8 => UNWINDOWED_710 ,
										MUX_10_1_IN_9 => UNWINDOWED_199 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_611
									);
MUX_REORD_UNIT_612 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_612 ,
										MUX_10_1_IN_1 => UNWINDOWED_612 ,
										MUX_10_1_IN_2 => UNWINDOWED_609 ,
										MUX_10_1_IN_3 => UNWINDOWED_616 ,
										MUX_10_1_IN_4 => UNWINDOWED_616 ,
										MUX_10_1_IN_5 => UNWINDOWED_585 ,
										MUX_10_1_IN_6 => UNWINDOWED_585 ,
										MUX_10_1_IN_7 => UNWINDOWED_712 ,
										MUX_10_1_IN_8 => UNWINDOWED_712 ,
										MUX_10_1_IN_9 => UNWINDOWED_201 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_612
									);
MUX_REORD_UNIT_613 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_613 ,
										MUX_10_1_IN_1 => UNWINDOWED_614 ,
										MUX_10_1_IN_2 => UNWINDOWED_611 ,
										MUX_10_1_IN_3 => UNWINDOWED_618 ,
										MUX_10_1_IN_4 => UNWINDOWED_618 ,
										MUX_10_1_IN_5 => UNWINDOWED_587 ,
										MUX_10_1_IN_6 => UNWINDOWED_587 ,
										MUX_10_1_IN_7 => UNWINDOWED_714 ,
										MUX_10_1_IN_8 => UNWINDOWED_714 ,
										MUX_10_1_IN_9 => UNWINDOWED_203 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_613
									);
MUX_REORD_UNIT_614 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_614 ,
										MUX_10_1_IN_1 => UNWINDOWED_613 ,
										MUX_10_1_IN_2 => UNWINDOWED_613 ,
										MUX_10_1_IN_3 => UNWINDOWED_620 ,
										MUX_10_1_IN_4 => UNWINDOWED_620 ,
										MUX_10_1_IN_5 => UNWINDOWED_589 ,
										MUX_10_1_IN_6 => UNWINDOWED_589 ,
										MUX_10_1_IN_7 => UNWINDOWED_716 ,
										MUX_10_1_IN_8 => UNWINDOWED_716 ,
										MUX_10_1_IN_9 => UNWINDOWED_205 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_614
									);
MUX_REORD_UNIT_615 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_615 ,
										MUX_10_1_IN_1 => UNWINDOWED_615 ,
										MUX_10_1_IN_2 => UNWINDOWED_615 ,
										MUX_10_1_IN_3 => UNWINDOWED_622 ,
										MUX_10_1_IN_4 => UNWINDOWED_622 ,
										MUX_10_1_IN_5 => UNWINDOWED_591 ,
										MUX_10_1_IN_6 => UNWINDOWED_591 ,
										MUX_10_1_IN_7 => UNWINDOWED_718 ,
										MUX_10_1_IN_8 => UNWINDOWED_718 ,
										MUX_10_1_IN_9 => UNWINDOWED_207 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_615
									);
MUX_REORD_UNIT_616 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_616 ,
										MUX_10_1_IN_1 => UNWINDOWED_616 ,
										MUX_10_1_IN_2 => UNWINDOWED_616 ,
										MUX_10_1_IN_3 => UNWINDOWED_609 ,
										MUX_10_1_IN_4 => UNWINDOWED_624 ,
										MUX_10_1_IN_5 => UNWINDOWED_593 ,
										MUX_10_1_IN_6 => UNWINDOWED_593 ,
										MUX_10_1_IN_7 => UNWINDOWED_720 ,
										MUX_10_1_IN_8 => UNWINDOWED_720 ,
										MUX_10_1_IN_9 => UNWINDOWED_209 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_616
									);
MUX_REORD_UNIT_617 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_617 ,
										MUX_10_1_IN_1 => UNWINDOWED_618 ,
										MUX_10_1_IN_2 => UNWINDOWED_618 ,
										MUX_10_1_IN_3 => UNWINDOWED_611 ,
										MUX_10_1_IN_4 => UNWINDOWED_626 ,
										MUX_10_1_IN_5 => UNWINDOWED_595 ,
										MUX_10_1_IN_6 => UNWINDOWED_595 ,
										MUX_10_1_IN_7 => UNWINDOWED_722 ,
										MUX_10_1_IN_8 => UNWINDOWED_722 ,
										MUX_10_1_IN_9 => UNWINDOWED_211 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_617
									);
MUX_REORD_UNIT_618 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_618 ,
										MUX_10_1_IN_1 => UNWINDOWED_617 ,
										MUX_10_1_IN_2 => UNWINDOWED_620 ,
										MUX_10_1_IN_3 => UNWINDOWED_613 ,
										MUX_10_1_IN_4 => UNWINDOWED_628 ,
										MUX_10_1_IN_5 => UNWINDOWED_597 ,
										MUX_10_1_IN_6 => UNWINDOWED_597 ,
										MUX_10_1_IN_7 => UNWINDOWED_724 ,
										MUX_10_1_IN_8 => UNWINDOWED_724 ,
										MUX_10_1_IN_9 => UNWINDOWED_213 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_618
									);
MUX_REORD_UNIT_619 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_619 ,
										MUX_10_1_IN_1 => UNWINDOWED_619 ,
										MUX_10_1_IN_2 => UNWINDOWED_622 ,
										MUX_10_1_IN_3 => UNWINDOWED_615 ,
										MUX_10_1_IN_4 => UNWINDOWED_630 ,
										MUX_10_1_IN_5 => UNWINDOWED_599 ,
										MUX_10_1_IN_6 => UNWINDOWED_599 ,
										MUX_10_1_IN_7 => UNWINDOWED_726 ,
										MUX_10_1_IN_8 => UNWINDOWED_726 ,
										MUX_10_1_IN_9 => UNWINDOWED_215 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_619
									);
MUX_REORD_UNIT_620 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_620 ,
										MUX_10_1_IN_1 => UNWINDOWED_620 ,
										MUX_10_1_IN_2 => UNWINDOWED_617 ,
										MUX_10_1_IN_3 => UNWINDOWED_617 ,
										MUX_10_1_IN_4 => UNWINDOWED_632 ,
										MUX_10_1_IN_5 => UNWINDOWED_601 ,
										MUX_10_1_IN_6 => UNWINDOWED_601 ,
										MUX_10_1_IN_7 => UNWINDOWED_728 ,
										MUX_10_1_IN_8 => UNWINDOWED_728 ,
										MUX_10_1_IN_9 => UNWINDOWED_217 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_620
									);
MUX_REORD_UNIT_621 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_621 ,
										MUX_10_1_IN_1 => UNWINDOWED_622 ,
										MUX_10_1_IN_2 => UNWINDOWED_619 ,
										MUX_10_1_IN_3 => UNWINDOWED_619 ,
										MUX_10_1_IN_4 => UNWINDOWED_634 ,
										MUX_10_1_IN_5 => UNWINDOWED_603 ,
										MUX_10_1_IN_6 => UNWINDOWED_603 ,
										MUX_10_1_IN_7 => UNWINDOWED_730 ,
										MUX_10_1_IN_8 => UNWINDOWED_730 ,
										MUX_10_1_IN_9 => UNWINDOWED_219 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_621
									);
MUX_REORD_UNIT_622 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_622 ,
										MUX_10_1_IN_1 => UNWINDOWED_621 ,
										MUX_10_1_IN_2 => UNWINDOWED_621 ,
										MUX_10_1_IN_3 => UNWINDOWED_621 ,
										MUX_10_1_IN_4 => UNWINDOWED_636 ,
										MUX_10_1_IN_5 => UNWINDOWED_605 ,
										MUX_10_1_IN_6 => UNWINDOWED_605 ,
										MUX_10_1_IN_7 => UNWINDOWED_732 ,
										MUX_10_1_IN_8 => UNWINDOWED_732 ,
										MUX_10_1_IN_9 => UNWINDOWED_221 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_622
									);
MUX_REORD_UNIT_623 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_623 ,
										MUX_10_1_IN_1 => UNWINDOWED_623 ,
										MUX_10_1_IN_2 => UNWINDOWED_623 ,
										MUX_10_1_IN_3 => UNWINDOWED_623 ,
										MUX_10_1_IN_4 => UNWINDOWED_638 ,
										MUX_10_1_IN_5 => UNWINDOWED_607 ,
										MUX_10_1_IN_6 => UNWINDOWED_607 ,
										MUX_10_1_IN_7 => UNWINDOWED_734 ,
										MUX_10_1_IN_8 => UNWINDOWED_734 ,
										MUX_10_1_IN_9 => UNWINDOWED_223 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_623
									);
MUX_REORD_UNIT_624 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_624 ,
										MUX_10_1_IN_1 => UNWINDOWED_624 ,
										MUX_10_1_IN_2 => UNWINDOWED_624 ,
										MUX_10_1_IN_3 => UNWINDOWED_624 ,
										MUX_10_1_IN_4 => UNWINDOWED_609 ,
										MUX_10_1_IN_5 => UNWINDOWED_609 ,
										MUX_10_1_IN_6 => UNWINDOWED_609 ,
										MUX_10_1_IN_7 => UNWINDOWED_736 ,
										MUX_10_1_IN_8 => UNWINDOWED_736 ,
										MUX_10_1_IN_9 => UNWINDOWED_225 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_624
									);
MUX_REORD_UNIT_625 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_625 ,
										MUX_10_1_IN_1 => UNWINDOWED_626 ,
										MUX_10_1_IN_2 => UNWINDOWED_626 ,
										MUX_10_1_IN_3 => UNWINDOWED_626 ,
										MUX_10_1_IN_4 => UNWINDOWED_611 ,
										MUX_10_1_IN_5 => UNWINDOWED_611 ,
										MUX_10_1_IN_6 => UNWINDOWED_611 ,
										MUX_10_1_IN_7 => UNWINDOWED_738 ,
										MUX_10_1_IN_8 => UNWINDOWED_738 ,
										MUX_10_1_IN_9 => UNWINDOWED_227 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_625
									);
MUX_REORD_UNIT_626 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_626 ,
										MUX_10_1_IN_1 => UNWINDOWED_625 ,
										MUX_10_1_IN_2 => UNWINDOWED_628 ,
										MUX_10_1_IN_3 => UNWINDOWED_628 ,
										MUX_10_1_IN_4 => UNWINDOWED_613 ,
										MUX_10_1_IN_5 => UNWINDOWED_613 ,
										MUX_10_1_IN_6 => UNWINDOWED_613 ,
										MUX_10_1_IN_7 => UNWINDOWED_740 ,
										MUX_10_1_IN_8 => UNWINDOWED_740 ,
										MUX_10_1_IN_9 => UNWINDOWED_229 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_626
									);
MUX_REORD_UNIT_627 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_627 ,
										MUX_10_1_IN_1 => UNWINDOWED_627 ,
										MUX_10_1_IN_2 => UNWINDOWED_630 ,
										MUX_10_1_IN_3 => UNWINDOWED_630 ,
										MUX_10_1_IN_4 => UNWINDOWED_615 ,
										MUX_10_1_IN_5 => UNWINDOWED_615 ,
										MUX_10_1_IN_6 => UNWINDOWED_615 ,
										MUX_10_1_IN_7 => UNWINDOWED_742 ,
										MUX_10_1_IN_8 => UNWINDOWED_742 ,
										MUX_10_1_IN_9 => UNWINDOWED_231 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_627
									);
MUX_REORD_UNIT_628 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_628 ,
										MUX_10_1_IN_1 => UNWINDOWED_628 ,
										MUX_10_1_IN_2 => UNWINDOWED_625 ,
										MUX_10_1_IN_3 => UNWINDOWED_632 ,
										MUX_10_1_IN_4 => UNWINDOWED_617 ,
										MUX_10_1_IN_5 => UNWINDOWED_617 ,
										MUX_10_1_IN_6 => UNWINDOWED_617 ,
										MUX_10_1_IN_7 => UNWINDOWED_744 ,
										MUX_10_1_IN_8 => UNWINDOWED_744 ,
										MUX_10_1_IN_9 => UNWINDOWED_233 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_628
									);
MUX_REORD_UNIT_629 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_629 ,
										MUX_10_1_IN_1 => UNWINDOWED_630 ,
										MUX_10_1_IN_2 => UNWINDOWED_627 ,
										MUX_10_1_IN_3 => UNWINDOWED_634 ,
										MUX_10_1_IN_4 => UNWINDOWED_619 ,
										MUX_10_1_IN_5 => UNWINDOWED_619 ,
										MUX_10_1_IN_6 => UNWINDOWED_619 ,
										MUX_10_1_IN_7 => UNWINDOWED_746 ,
										MUX_10_1_IN_8 => UNWINDOWED_746 ,
										MUX_10_1_IN_9 => UNWINDOWED_235 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_629
									);
MUX_REORD_UNIT_630 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_630 ,
										MUX_10_1_IN_1 => UNWINDOWED_629 ,
										MUX_10_1_IN_2 => UNWINDOWED_629 ,
										MUX_10_1_IN_3 => UNWINDOWED_636 ,
										MUX_10_1_IN_4 => UNWINDOWED_621 ,
										MUX_10_1_IN_5 => UNWINDOWED_621 ,
										MUX_10_1_IN_6 => UNWINDOWED_621 ,
										MUX_10_1_IN_7 => UNWINDOWED_748 ,
										MUX_10_1_IN_8 => UNWINDOWED_748 ,
										MUX_10_1_IN_9 => UNWINDOWED_237 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_630
									);
MUX_REORD_UNIT_631 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_631 ,
										MUX_10_1_IN_1 => UNWINDOWED_631 ,
										MUX_10_1_IN_2 => UNWINDOWED_631 ,
										MUX_10_1_IN_3 => UNWINDOWED_638 ,
										MUX_10_1_IN_4 => UNWINDOWED_623 ,
										MUX_10_1_IN_5 => UNWINDOWED_623 ,
										MUX_10_1_IN_6 => UNWINDOWED_623 ,
										MUX_10_1_IN_7 => UNWINDOWED_750 ,
										MUX_10_1_IN_8 => UNWINDOWED_750 ,
										MUX_10_1_IN_9 => UNWINDOWED_239 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_631
									);
MUX_REORD_UNIT_632 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_632 ,
										MUX_10_1_IN_1 => UNWINDOWED_632 ,
										MUX_10_1_IN_2 => UNWINDOWED_632 ,
										MUX_10_1_IN_3 => UNWINDOWED_625 ,
										MUX_10_1_IN_4 => UNWINDOWED_625 ,
										MUX_10_1_IN_5 => UNWINDOWED_625 ,
										MUX_10_1_IN_6 => UNWINDOWED_625 ,
										MUX_10_1_IN_7 => UNWINDOWED_752 ,
										MUX_10_1_IN_8 => UNWINDOWED_752 ,
										MUX_10_1_IN_9 => UNWINDOWED_241 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_632
									);
MUX_REORD_UNIT_633 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_633 ,
										MUX_10_1_IN_1 => UNWINDOWED_634 ,
										MUX_10_1_IN_2 => UNWINDOWED_634 ,
										MUX_10_1_IN_3 => UNWINDOWED_627 ,
										MUX_10_1_IN_4 => UNWINDOWED_627 ,
										MUX_10_1_IN_5 => UNWINDOWED_627 ,
										MUX_10_1_IN_6 => UNWINDOWED_627 ,
										MUX_10_1_IN_7 => UNWINDOWED_754 ,
										MUX_10_1_IN_8 => UNWINDOWED_754 ,
										MUX_10_1_IN_9 => UNWINDOWED_243 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_633
									);
MUX_REORD_UNIT_634 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_634 ,
										MUX_10_1_IN_1 => UNWINDOWED_633 ,
										MUX_10_1_IN_2 => UNWINDOWED_636 ,
										MUX_10_1_IN_3 => UNWINDOWED_629 ,
										MUX_10_1_IN_4 => UNWINDOWED_629 ,
										MUX_10_1_IN_5 => UNWINDOWED_629 ,
										MUX_10_1_IN_6 => UNWINDOWED_629 ,
										MUX_10_1_IN_7 => UNWINDOWED_756 ,
										MUX_10_1_IN_8 => UNWINDOWED_756 ,
										MUX_10_1_IN_9 => UNWINDOWED_245 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_634
									);
MUX_REORD_UNIT_635 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_635 ,
										MUX_10_1_IN_1 => UNWINDOWED_635 ,
										MUX_10_1_IN_2 => UNWINDOWED_638 ,
										MUX_10_1_IN_3 => UNWINDOWED_631 ,
										MUX_10_1_IN_4 => UNWINDOWED_631 ,
										MUX_10_1_IN_5 => UNWINDOWED_631 ,
										MUX_10_1_IN_6 => UNWINDOWED_631 ,
										MUX_10_1_IN_7 => UNWINDOWED_758 ,
										MUX_10_1_IN_8 => UNWINDOWED_758 ,
										MUX_10_1_IN_9 => UNWINDOWED_247 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_635
									);
MUX_REORD_UNIT_636 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_636 ,
										MUX_10_1_IN_1 => UNWINDOWED_636 ,
										MUX_10_1_IN_2 => UNWINDOWED_633 ,
										MUX_10_1_IN_3 => UNWINDOWED_633 ,
										MUX_10_1_IN_4 => UNWINDOWED_633 ,
										MUX_10_1_IN_5 => UNWINDOWED_633 ,
										MUX_10_1_IN_6 => UNWINDOWED_633 ,
										MUX_10_1_IN_7 => UNWINDOWED_760 ,
										MUX_10_1_IN_8 => UNWINDOWED_760 ,
										MUX_10_1_IN_9 => UNWINDOWED_249 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_636
									);
MUX_REORD_UNIT_637 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_637 ,
										MUX_10_1_IN_1 => UNWINDOWED_638 ,
										MUX_10_1_IN_2 => UNWINDOWED_635 ,
										MUX_10_1_IN_3 => UNWINDOWED_635 ,
										MUX_10_1_IN_4 => UNWINDOWED_635 ,
										MUX_10_1_IN_5 => UNWINDOWED_635 ,
										MUX_10_1_IN_6 => UNWINDOWED_635 ,
										MUX_10_1_IN_7 => UNWINDOWED_762 ,
										MUX_10_1_IN_8 => UNWINDOWED_762 ,
										MUX_10_1_IN_9 => UNWINDOWED_251 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_637
									);
MUX_REORD_UNIT_638 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_638 ,
										MUX_10_1_IN_1 => UNWINDOWED_637 ,
										MUX_10_1_IN_2 => UNWINDOWED_637 ,
										MUX_10_1_IN_3 => UNWINDOWED_637 ,
										MUX_10_1_IN_4 => UNWINDOWED_637 ,
										MUX_10_1_IN_5 => UNWINDOWED_637 ,
										MUX_10_1_IN_6 => UNWINDOWED_637 ,
										MUX_10_1_IN_7 => UNWINDOWED_764 ,
										MUX_10_1_IN_8 => UNWINDOWED_764 ,
										MUX_10_1_IN_9 => UNWINDOWED_253 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_638
									);
MUX_REORD_UNIT_639 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_639 ,
										MUX_10_1_IN_1 => UNWINDOWED_639 ,
										MUX_10_1_IN_2 => UNWINDOWED_639 ,
										MUX_10_1_IN_3 => UNWINDOWED_639 ,
										MUX_10_1_IN_4 => UNWINDOWED_639 ,
										MUX_10_1_IN_5 => UNWINDOWED_639 ,
										MUX_10_1_IN_6 => UNWINDOWED_639 ,
										MUX_10_1_IN_7 => UNWINDOWED_766 ,
										MUX_10_1_IN_8 => UNWINDOWED_766 ,
										MUX_10_1_IN_9 => UNWINDOWED_255 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_639
									);
MUX_REORD_UNIT_640 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_640 ,
										MUX_10_1_IN_1 => UNWINDOWED_640 ,
										MUX_10_1_IN_2 => UNWINDOWED_640 ,
										MUX_10_1_IN_3 => UNWINDOWED_640 ,
										MUX_10_1_IN_4 => UNWINDOWED_640 ,
										MUX_10_1_IN_5 => UNWINDOWED_640 ,
										MUX_10_1_IN_6 => UNWINDOWED_640 ,
										MUX_10_1_IN_7 => UNWINDOWED_513 ,
										MUX_10_1_IN_8 => UNWINDOWED_768 ,
										MUX_10_1_IN_9 => UNWINDOWED_257 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_640
									);
MUX_REORD_UNIT_641 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_641 ,
										MUX_10_1_IN_1 => UNWINDOWED_642 ,
										MUX_10_1_IN_2 => UNWINDOWED_642 ,
										MUX_10_1_IN_3 => UNWINDOWED_642 ,
										MUX_10_1_IN_4 => UNWINDOWED_642 ,
										MUX_10_1_IN_5 => UNWINDOWED_642 ,
										MUX_10_1_IN_6 => UNWINDOWED_642 ,
										MUX_10_1_IN_7 => UNWINDOWED_515 ,
										MUX_10_1_IN_8 => UNWINDOWED_770 ,
										MUX_10_1_IN_9 => UNWINDOWED_259 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_641
									);
MUX_REORD_UNIT_642 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_642 ,
										MUX_10_1_IN_1 => UNWINDOWED_641 ,
										MUX_10_1_IN_2 => UNWINDOWED_644 ,
										MUX_10_1_IN_3 => UNWINDOWED_644 ,
										MUX_10_1_IN_4 => UNWINDOWED_644 ,
										MUX_10_1_IN_5 => UNWINDOWED_644 ,
										MUX_10_1_IN_6 => UNWINDOWED_644 ,
										MUX_10_1_IN_7 => UNWINDOWED_517 ,
										MUX_10_1_IN_8 => UNWINDOWED_772 ,
										MUX_10_1_IN_9 => UNWINDOWED_261 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_642
									);
MUX_REORD_UNIT_643 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_643 ,
										MUX_10_1_IN_1 => UNWINDOWED_643 ,
										MUX_10_1_IN_2 => UNWINDOWED_646 ,
										MUX_10_1_IN_3 => UNWINDOWED_646 ,
										MUX_10_1_IN_4 => UNWINDOWED_646 ,
										MUX_10_1_IN_5 => UNWINDOWED_646 ,
										MUX_10_1_IN_6 => UNWINDOWED_646 ,
										MUX_10_1_IN_7 => UNWINDOWED_519 ,
										MUX_10_1_IN_8 => UNWINDOWED_774 ,
										MUX_10_1_IN_9 => UNWINDOWED_263 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_643
									);
MUX_REORD_UNIT_644 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_644 ,
										MUX_10_1_IN_1 => UNWINDOWED_644 ,
										MUX_10_1_IN_2 => UNWINDOWED_641 ,
										MUX_10_1_IN_3 => UNWINDOWED_648 ,
										MUX_10_1_IN_4 => UNWINDOWED_648 ,
										MUX_10_1_IN_5 => UNWINDOWED_648 ,
										MUX_10_1_IN_6 => UNWINDOWED_648 ,
										MUX_10_1_IN_7 => UNWINDOWED_521 ,
										MUX_10_1_IN_8 => UNWINDOWED_776 ,
										MUX_10_1_IN_9 => UNWINDOWED_265 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_644
									);
MUX_REORD_UNIT_645 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_645 ,
										MUX_10_1_IN_1 => UNWINDOWED_646 ,
										MUX_10_1_IN_2 => UNWINDOWED_643 ,
										MUX_10_1_IN_3 => UNWINDOWED_650 ,
										MUX_10_1_IN_4 => UNWINDOWED_650 ,
										MUX_10_1_IN_5 => UNWINDOWED_650 ,
										MUX_10_1_IN_6 => UNWINDOWED_650 ,
										MUX_10_1_IN_7 => UNWINDOWED_523 ,
										MUX_10_1_IN_8 => UNWINDOWED_778 ,
										MUX_10_1_IN_9 => UNWINDOWED_267 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_645
									);
MUX_REORD_UNIT_646 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_646 ,
										MUX_10_1_IN_1 => UNWINDOWED_645 ,
										MUX_10_1_IN_2 => UNWINDOWED_645 ,
										MUX_10_1_IN_3 => UNWINDOWED_652 ,
										MUX_10_1_IN_4 => UNWINDOWED_652 ,
										MUX_10_1_IN_5 => UNWINDOWED_652 ,
										MUX_10_1_IN_6 => UNWINDOWED_652 ,
										MUX_10_1_IN_7 => UNWINDOWED_525 ,
										MUX_10_1_IN_8 => UNWINDOWED_780 ,
										MUX_10_1_IN_9 => UNWINDOWED_269 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_646
									);
MUX_REORD_UNIT_647 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_647 ,
										MUX_10_1_IN_1 => UNWINDOWED_647 ,
										MUX_10_1_IN_2 => UNWINDOWED_647 ,
										MUX_10_1_IN_3 => UNWINDOWED_654 ,
										MUX_10_1_IN_4 => UNWINDOWED_654 ,
										MUX_10_1_IN_5 => UNWINDOWED_654 ,
										MUX_10_1_IN_6 => UNWINDOWED_654 ,
										MUX_10_1_IN_7 => UNWINDOWED_527 ,
										MUX_10_1_IN_8 => UNWINDOWED_782 ,
										MUX_10_1_IN_9 => UNWINDOWED_271 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_647
									);
MUX_REORD_UNIT_648 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_648 ,
										MUX_10_1_IN_1 => UNWINDOWED_648 ,
										MUX_10_1_IN_2 => UNWINDOWED_648 ,
										MUX_10_1_IN_3 => UNWINDOWED_641 ,
										MUX_10_1_IN_4 => UNWINDOWED_656 ,
										MUX_10_1_IN_5 => UNWINDOWED_656 ,
										MUX_10_1_IN_6 => UNWINDOWED_656 ,
										MUX_10_1_IN_7 => UNWINDOWED_529 ,
										MUX_10_1_IN_8 => UNWINDOWED_784 ,
										MUX_10_1_IN_9 => UNWINDOWED_273 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_648
									);
MUX_REORD_UNIT_649 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_649 ,
										MUX_10_1_IN_1 => UNWINDOWED_650 ,
										MUX_10_1_IN_2 => UNWINDOWED_650 ,
										MUX_10_1_IN_3 => UNWINDOWED_643 ,
										MUX_10_1_IN_4 => UNWINDOWED_658 ,
										MUX_10_1_IN_5 => UNWINDOWED_658 ,
										MUX_10_1_IN_6 => UNWINDOWED_658 ,
										MUX_10_1_IN_7 => UNWINDOWED_531 ,
										MUX_10_1_IN_8 => UNWINDOWED_786 ,
										MUX_10_1_IN_9 => UNWINDOWED_275 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_649
									);
MUX_REORD_UNIT_650 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_650 ,
										MUX_10_1_IN_1 => UNWINDOWED_649 ,
										MUX_10_1_IN_2 => UNWINDOWED_652 ,
										MUX_10_1_IN_3 => UNWINDOWED_645 ,
										MUX_10_1_IN_4 => UNWINDOWED_660 ,
										MUX_10_1_IN_5 => UNWINDOWED_660 ,
										MUX_10_1_IN_6 => UNWINDOWED_660 ,
										MUX_10_1_IN_7 => UNWINDOWED_533 ,
										MUX_10_1_IN_8 => UNWINDOWED_788 ,
										MUX_10_1_IN_9 => UNWINDOWED_277 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_650
									);
MUX_REORD_UNIT_651 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_651 ,
										MUX_10_1_IN_1 => UNWINDOWED_651 ,
										MUX_10_1_IN_2 => UNWINDOWED_654 ,
										MUX_10_1_IN_3 => UNWINDOWED_647 ,
										MUX_10_1_IN_4 => UNWINDOWED_662 ,
										MUX_10_1_IN_5 => UNWINDOWED_662 ,
										MUX_10_1_IN_6 => UNWINDOWED_662 ,
										MUX_10_1_IN_7 => UNWINDOWED_535 ,
										MUX_10_1_IN_8 => UNWINDOWED_790 ,
										MUX_10_1_IN_9 => UNWINDOWED_279 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_651
									);
MUX_REORD_UNIT_652 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_652 ,
										MUX_10_1_IN_1 => UNWINDOWED_652 ,
										MUX_10_1_IN_2 => UNWINDOWED_649 ,
										MUX_10_1_IN_3 => UNWINDOWED_649 ,
										MUX_10_1_IN_4 => UNWINDOWED_664 ,
										MUX_10_1_IN_5 => UNWINDOWED_664 ,
										MUX_10_1_IN_6 => UNWINDOWED_664 ,
										MUX_10_1_IN_7 => UNWINDOWED_537 ,
										MUX_10_1_IN_8 => UNWINDOWED_792 ,
										MUX_10_1_IN_9 => UNWINDOWED_281 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_652
									);
MUX_REORD_UNIT_653 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_653 ,
										MUX_10_1_IN_1 => UNWINDOWED_654 ,
										MUX_10_1_IN_2 => UNWINDOWED_651 ,
										MUX_10_1_IN_3 => UNWINDOWED_651 ,
										MUX_10_1_IN_4 => UNWINDOWED_666 ,
										MUX_10_1_IN_5 => UNWINDOWED_666 ,
										MUX_10_1_IN_6 => UNWINDOWED_666 ,
										MUX_10_1_IN_7 => UNWINDOWED_539 ,
										MUX_10_1_IN_8 => UNWINDOWED_794 ,
										MUX_10_1_IN_9 => UNWINDOWED_283 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_653
									);
MUX_REORD_UNIT_654 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_654 ,
										MUX_10_1_IN_1 => UNWINDOWED_653 ,
										MUX_10_1_IN_2 => UNWINDOWED_653 ,
										MUX_10_1_IN_3 => UNWINDOWED_653 ,
										MUX_10_1_IN_4 => UNWINDOWED_668 ,
										MUX_10_1_IN_5 => UNWINDOWED_668 ,
										MUX_10_1_IN_6 => UNWINDOWED_668 ,
										MUX_10_1_IN_7 => UNWINDOWED_541 ,
										MUX_10_1_IN_8 => UNWINDOWED_796 ,
										MUX_10_1_IN_9 => UNWINDOWED_285 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_654
									);
MUX_REORD_UNIT_655 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_655 ,
										MUX_10_1_IN_1 => UNWINDOWED_655 ,
										MUX_10_1_IN_2 => UNWINDOWED_655 ,
										MUX_10_1_IN_3 => UNWINDOWED_655 ,
										MUX_10_1_IN_4 => UNWINDOWED_670 ,
										MUX_10_1_IN_5 => UNWINDOWED_670 ,
										MUX_10_1_IN_6 => UNWINDOWED_670 ,
										MUX_10_1_IN_7 => UNWINDOWED_543 ,
										MUX_10_1_IN_8 => UNWINDOWED_798 ,
										MUX_10_1_IN_9 => UNWINDOWED_287 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_655
									);
MUX_REORD_UNIT_656 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_656 ,
										MUX_10_1_IN_1 => UNWINDOWED_656 ,
										MUX_10_1_IN_2 => UNWINDOWED_656 ,
										MUX_10_1_IN_3 => UNWINDOWED_656 ,
										MUX_10_1_IN_4 => UNWINDOWED_641 ,
										MUX_10_1_IN_5 => UNWINDOWED_672 ,
										MUX_10_1_IN_6 => UNWINDOWED_672 ,
										MUX_10_1_IN_7 => UNWINDOWED_545 ,
										MUX_10_1_IN_8 => UNWINDOWED_800 ,
										MUX_10_1_IN_9 => UNWINDOWED_289 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_656
									);
MUX_REORD_UNIT_657 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_657 ,
										MUX_10_1_IN_1 => UNWINDOWED_658 ,
										MUX_10_1_IN_2 => UNWINDOWED_658 ,
										MUX_10_1_IN_3 => UNWINDOWED_658 ,
										MUX_10_1_IN_4 => UNWINDOWED_643 ,
										MUX_10_1_IN_5 => UNWINDOWED_674 ,
										MUX_10_1_IN_6 => UNWINDOWED_674 ,
										MUX_10_1_IN_7 => UNWINDOWED_547 ,
										MUX_10_1_IN_8 => UNWINDOWED_802 ,
										MUX_10_1_IN_9 => UNWINDOWED_291 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_657
									);
MUX_REORD_UNIT_658 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_658 ,
										MUX_10_1_IN_1 => UNWINDOWED_657 ,
										MUX_10_1_IN_2 => UNWINDOWED_660 ,
										MUX_10_1_IN_3 => UNWINDOWED_660 ,
										MUX_10_1_IN_4 => UNWINDOWED_645 ,
										MUX_10_1_IN_5 => UNWINDOWED_676 ,
										MUX_10_1_IN_6 => UNWINDOWED_676 ,
										MUX_10_1_IN_7 => UNWINDOWED_549 ,
										MUX_10_1_IN_8 => UNWINDOWED_804 ,
										MUX_10_1_IN_9 => UNWINDOWED_293 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_658
									);
MUX_REORD_UNIT_659 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_659 ,
										MUX_10_1_IN_1 => UNWINDOWED_659 ,
										MUX_10_1_IN_2 => UNWINDOWED_662 ,
										MUX_10_1_IN_3 => UNWINDOWED_662 ,
										MUX_10_1_IN_4 => UNWINDOWED_647 ,
										MUX_10_1_IN_5 => UNWINDOWED_678 ,
										MUX_10_1_IN_6 => UNWINDOWED_678 ,
										MUX_10_1_IN_7 => UNWINDOWED_551 ,
										MUX_10_1_IN_8 => UNWINDOWED_806 ,
										MUX_10_1_IN_9 => UNWINDOWED_295 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_659
									);
MUX_REORD_UNIT_660 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_660 ,
										MUX_10_1_IN_1 => UNWINDOWED_660 ,
										MUX_10_1_IN_2 => UNWINDOWED_657 ,
										MUX_10_1_IN_3 => UNWINDOWED_664 ,
										MUX_10_1_IN_4 => UNWINDOWED_649 ,
										MUX_10_1_IN_5 => UNWINDOWED_680 ,
										MUX_10_1_IN_6 => UNWINDOWED_680 ,
										MUX_10_1_IN_7 => UNWINDOWED_553 ,
										MUX_10_1_IN_8 => UNWINDOWED_808 ,
										MUX_10_1_IN_9 => UNWINDOWED_297 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_660
									);
MUX_REORD_UNIT_661 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_661 ,
										MUX_10_1_IN_1 => UNWINDOWED_662 ,
										MUX_10_1_IN_2 => UNWINDOWED_659 ,
										MUX_10_1_IN_3 => UNWINDOWED_666 ,
										MUX_10_1_IN_4 => UNWINDOWED_651 ,
										MUX_10_1_IN_5 => UNWINDOWED_682 ,
										MUX_10_1_IN_6 => UNWINDOWED_682 ,
										MUX_10_1_IN_7 => UNWINDOWED_555 ,
										MUX_10_1_IN_8 => UNWINDOWED_810 ,
										MUX_10_1_IN_9 => UNWINDOWED_299 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_661
									);
MUX_REORD_UNIT_662 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_662 ,
										MUX_10_1_IN_1 => UNWINDOWED_661 ,
										MUX_10_1_IN_2 => UNWINDOWED_661 ,
										MUX_10_1_IN_3 => UNWINDOWED_668 ,
										MUX_10_1_IN_4 => UNWINDOWED_653 ,
										MUX_10_1_IN_5 => UNWINDOWED_684 ,
										MUX_10_1_IN_6 => UNWINDOWED_684 ,
										MUX_10_1_IN_7 => UNWINDOWED_557 ,
										MUX_10_1_IN_8 => UNWINDOWED_812 ,
										MUX_10_1_IN_9 => UNWINDOWED_301 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_662
									);
MUX_REORD_UNIT_663 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_663 ,
										MUX_10_1_IN_1 => UNWINDOWED_663 ,
										MUX_10_1_IN_2 => UNWINDOWED_663 ,
										MUX_10_1_IN_3 => UNWINDOWED_670 ,
										MUX_10_1_IN_4 => UNWINDOWED_655 ,
										MUX_10_1_IN_5 => UNWINDOWED_686 ,
										MUX_10_1_IN_6 => UNWINDOWED_686 ,
										MUX_10_1_IN_7 => UNWINDOWED_559 ,
										MUX_10_1_IN_8 => UNWINDOWED_814 ,
										MUX_10_1_IN_9 => UNWINDOWED_303 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_663
									);
MUX_REORD_UNIT_664 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_664 ,
										MUX_10_1_IN_1 => UNWINDOWED_664 ,
										MUX_10_1_IN_2 => UNWINDOWED_664 ,
										MUX_10_1_IN_3 => UNWINDOWED_657 ,
										MUX_10_1_IN_4 => UNWINDOWED_657 ,
										MUX_10_1_IN_5 => UNWINDOWED_688 ,
										MUX_10_1_IN_6 => UNWINDOWED_688 ,
										MUX_10_1_IN_7 => UNWINDOWED_561 ,
										MUX_10_1_IN_8 => UNWINDOWED_816 ,
										MUX_10_1_IN_9 => UNWINDOWED_305 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_664
									);
MUX_REORD_UNIT_665 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_665 ,
										MUX_10_1_IN_1 => UNWINDOWED_666 ,
										MUX_10_1_IN_2 => UNWINDOWED_666 ,
										MUX_10_1_IN_3 => UNWINDOWED_659 ,
										MUX_10_1_IN_4 => UNWINDOWED_659 ,
										MUX_10_1_IN_5 => UNWINDOWED_690 ,
										MUX_10_1_IN_6 => UNWINDOWED_690 ,
										MUX_10_1_IN_7 => UNWINDOWED_563 ,
										MUX_10_1_IN_8 => UNWINDOWED_818 ,
										MUX_10_1_IN_9 => UNWINDOWED_307 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_665
									);
MUX_REORD_UNIT_666 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_666 ,
										MUX_10_1_IN_1 => UNWINDOWED_665 ,
										MUX_10_1_IN_2 => UNWINDOWED_668 ,
										MUX_10_1_IN_3 => UNWINDOWED_661 ,
										MUX_10_1_IN_4 => UNWINDOWED_661 ,
										MUX_10_1_IN_5 => UNWINDOWED_692 ,
										MUX_10_1_IN_6 => UNWINDOWED_692 ,
										MUX_10_1_IN_7 => UNWINDOWED_565 ,
										MUX_10_1_IN_8 => UNWINDOWED_820 ,
										MUX_10_1_IN_9 => UNWINDOWED_309 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_666
									);
MUX_REORD_UNIT_667 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_667 ,
										MUX_10_1_IN_1 => UNWINDOWED_667 ,
										MUX_10_1_IN_2 => UNWINDOWED_670 ,
										MUX_10_1_IN_3 => UNWINDOWED_663 ,
										MUX_10_1_IN_4 => UNWINDOWED_663 ,
										MUX_10_1_IN_5 => UNWINDOWED_694 ,
										MUX_10_1_IN_6 => UNWINDOWED_694 ,
										MUX_10_1_IN_7 => UNWINDOWED_567 ,
										MUX_10_1_IN_8 => UNWINDOWED_822 ,
										MUX_10_1_IN_9 => UNWINDOWED_311 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_667
									);
MUX_REORD_UNIT_668 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_668 ,
										MUX_10_1_IN_1 => UNWINDOWED_668 ,
										MUX_10_1_IN_2 => UNWINDOWED_665 ,
										MUX_10_1_IN_3 => UNWINDOWED_665 ,
										MUX_10_1_IN_4 => UNWINDOWED_665 ,
										MUX_10_1_IN_5 => UNWINDOWED_696 ,
										MUX_10_1_IN_6 => UNWINDOWED_696 ,
										MUX_10_1_IN_7 => UNWINDOWED_569 ,
										MUX_10_1_IN_8 => UNWINDOWED_824 ,
										MUX_10_1_IN_9 => UNWINDOWED_313 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_668
									);
MUX_REORD_UNIT_669 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_669 ,
										MUX_10_1_IN_1 => UNWINDOWED_670 ,
										MUX_10_1_IN_2 => UNWINDOWED_667 ,
										MUX_10_1_IN_3 => UNWINDOWED_667 ,
										MUX_10_1_IN_4 => UNWINDOWED_667 ,
										MUX_10_1_IN_5 => UNWINDOWED_698 ,
										MUX_10_1_IN_6 => UNWINDOWED_698 ,
										MUX_10_1_IN_7 => UNWINDOWED_571 ,
										MUX_10_1_IN_8 => UNWINDOWED_826 ,
										MUX_10_1_IN_9 => UNWINDOWED_315 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_669
									);
MUX_REORD_UNIT_670 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_670 ,
										MUX_10_1_IN_1 => UNWINDOWED_669 ,
										MUX_10_1_IN_2 => UNWINDOWED_669 ,
										MUX_10_1_IN_3 => UNWINDOWED_669 ,
										MUX_10_1_IN_4 => UNWINDOWED_669 ,
										MUX_10_1_IN_5 => UNWINDOWED_700 ,
										MUX_10_1_IN_6 => UNWINDOWED_700 ,
										MUX_10_1_IN_7 => UNWINDOWED_573 ,
										MUX_10_1_IN_8 => UNWINDOWED_828 ,
										MUX_10_1_IN_9 => UNWINDOWED_317 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_670
									);
MUX_REORD_UNIT_671 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_671 ,
										MUX_10_1_IN_1 => UNWINDOWED_671 ,
										MUX_10_1_IN_2 => UNWINDOWED_671 ,
										MUX_10_1_IN_3 => UNWINDOWED_671 ,
										MUX_10_1_IN_4 => UNWINDOWED_671 ,
										MUX_10_1_IN_5 => UNWINDOWED_702 ,
										MUX_10_1_IN_6 => UNWINDOWED_702 ,
										MUX_10_1_IN_7 => UNWINDOWED_575 ,
										MUX_10_1_IN_8 => UNWINDOWED_830 ,
										MUX_10_1_IN_9 => UNWINDOWED_319 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_671
									);
MUX_REORD_UNIT_672 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_672 ,
										MUX_10_1_IN_1 => UNWINDOWED_672 ,
										MUX_10_1_IN_2 => UNWINDOWED_672 ,
										MUX_10_1_IN_3 => UNWINDOWED_672 ,
										MUX_10_1_IN_4 => UNWINDOWED_672 ,
										MUX_10_1_IN_5 => UNWINDOWED_641 ,
										MUX_10_1_IN_6 => UNWINDOWED_704 ,
										MUX_10_1_IN_7 => UNWINDOWED_577 ,
										MUX_10_1_IN_8 => UNWINDOWED_832 ,
										MUX_10_1_IN_9 => UNWINDOWED_321 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_672
									);
MUX_REORD_UNIT_673 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_673 ,
										MUX_10_1_IN_1 => UNWINDOWED_674 ,
										MUX_10_1_IN_2 => UNWINDOWED_674 ,
										MUX_10_1_IN_3 => UNWINDOWED_674 ,
										MUX_10_1_IN_4 => UNWINDOWED_674 ,
										MUX_10_1_IN_5 => UNWINDOWED_643 ,
										MUX_10_1_IN_6 => UNWINDOWED_706 ,
										MUX_10_1_IN_7 => UNWINDOWED_579 ,
										MUX_10_1_IN_8 => UNWINDOWED_834 ,
										MUX_10_1_IN_9 => UNWINDOWED_323 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_673
									);
MUX_REORD_UNIT_674 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_674 ,
										MUX_10_1_IN_1 => UNWINDOWED_673 ,
										MUX_10_1_IN_2 => UNWINDOWED_676 ,
										MUX_10_1_IN_3 => UNWINDOWED_676 ,
										MUX_10_1_IN_4 => UNWINDOWED_676 ,
										MUX_10_1_IN_5 => UNWINDOWED_645 ,
										MUX_10_1_IN_6 => UNWINDOWED_708 ,
										MUX_10_1_IN_7 => UNWINDOWED_581 ,
										MUX_10_1_IN_8 => UNWINDOWED_836 ,
										MUX_10_1_IN_9 => UNWINDOWED_325 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_674
									);
MUX_REORD_UNIT_675 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_675 ,
										MUX_10_1_IN_1 => UNWINDOWED_675 ,
										MUX_10_1_IN_2 => UNWINDOWED_678 ,
										MUX_10_1_IN_3 => UNWINDOWED_678 ,
										MUX_10_1_IN_4 => UNWINDOWED_678 ,
										MUX_10_1_IN_5 => UNWINDOWED_647 ,
										MUX_10_1_IN_6 => UNWINDOWED_710 ,
										MUX_10_1_IN_7 => UNWINDOWED_583 ,
										MUX_10_1_IN_8 => UNWINDOWED_838 ,
										MUX_10_1_IN_9 => UNWINDOWED_327 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_675
									);
MUX_REORD_UNIT_676 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_676 ,
										MUX_10_1_IN_1 => UNWINDOWED_676 ,
										MUX_10_1_IN_2 => UNWINDOWED_673 ,
										MUX_10_1_IN_3 => UNWINDOWED_680 ,
										MUX_10_1_IN_4 => UNWINDOWED_680 ,
										MUX_10_1_IN_5 => UNWINDOWED_649 ,
										MUX_10_1_IN_6 => UNWINDOWED_712 ,
										MUX_10_1_IN_7 => UNWINDOWED_585 ,
										MUX_10_1_IN_8 => UNWINDOWED_840 ,
										MUX_10_1_IN_9 => UNWINDOWED_329 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_676
									);
MUX_REORD_UNIT_677 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_677 ,
										MUX_10_1_IN_1 => UNWINDOWED_678 ,
										MUX_10_1_IN_2 => UNWINDOWED_675 ,
										MUX_10_1_IN_3 => UNWINDOWED_682 ,
										MUX_10_1_IN_4 => UNWINDOWED_682 ,
										MUX_10_1_IN_5 => UNWINDOWED_651 ,
										MUX_10_1_IN_6 => UNWINDOWED_714 ,
										MUX_10_1_IN_7 => UNWINDOWED_587 ,
										MUX_10_1_IN_8 => UNWINDOWED_842 ,
										MUX_10_1_IN_9 => UNWINDOWED_331 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_677
									);
MUX_REORD_UNIT_678 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_678 ,
										MUX_10_1_IN_1 => UNWINDOWED_677 ,
										MUX_10_1_IN_2 => UNWINDOWED_677 ,
										MUX_10_1_IN_3 => UNWINDOWED_684 ,
										MUX_10_1_IN_4 => UNWINDOWED_684 ,
										MUX_10_1_IN_5 => UNWINDOWED_653 ,
										MUX_10_1_IN_6 => UNWINDOWED_716 ,
										MUX_10_1_IN_7 => UNWINDOWED_589 ,
										MUX_10_1_IN_8 => UNWINDOWED_844 ,
										MUX_10_1_IN_9 => UNWINDOWED_333 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_678
									);
MUX_REORD_UNIT_679 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_679 ,
										MUX_10_1_IN_1 => UNWINDOWED_679 ,
										MUX_10_1_IN_2 => UNWINDOWED_679 ,
										MUX_10_1_IN_3 => UNWINDOWED_686 ,
										MUX_10_1_IN_4 => UNWINDOWED_686 ,
										MUX_10_1_IN_5 => UNWINDOWED_655 ,
										MUX_10_1_IN_6 => UNWINDOWED_718 ,
										MUX_10_1_IN_7 => UNWINDOWED_591 ,
										MUX_10_1_IN_8 => UNWINDOWED_846 ,
										MUX_10_1_IN_9 => UNWINDOWED_335 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_679
									);
MUX_REORD_UNIT_680 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_680 ,
										MUX_10_1_IN_1 => UNWINDOWED_680 ,
										MUX_10_1_IN_2 => UNWINDOWED_680 ,
										MUX_10_1_IN_3 => UNWINDOWED_673 ,
										MUX_10_1_IN_4 => UNWINDOWED_688 ,
										MUX_10_1_IN_5 => UNWINDOWED_657 ,
										MUX_10_1_IN_6 => UNWINDOWED_720 ,
										MUX_10_1_IN_7 => UNWINDOWED_593 ,
										MUX_10_1_IN_8 => UNWINDOWED_848 ,
										MUX_10_1_IN_9 => UNWINDOWED_337 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_680
									);
MUX_REORD_UNIT_681 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_681 ,
										MUX_10_1_IN_1 => UNWINDOWED_682 ,
										MUX_10_1_IN_2 => UNWINDOWED_682 ,
										MUX_10_1_IN_3 => UNWINDOWED_675 ,
										MUX_10_1_IN_4 => UNWINDOWED_690 ,
										MUX_10_1_IN_5 => UNWINDOWED_659 ,
										MUX_10_1_IN_6 => UNWINDOWED_722 ,
										MUX_10_1_IN_7 => UNWINDOWED_595 ,
										MUX_10_1_IN_8 => UNWINDOWED_850 ,
										MUX_10_1_IN_9 => UNWINDOWED_339 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_681
									);
MUX_REORD_UNIT_682 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_682 ,
										MUX_10_1_IN_1 => UNWINDOWED_681 ,
										MUX_10_1_IN_2 => UNWINDOWED_684 ,
										MUX_10_1_IN_3 => UNWINDOWED_677 ,
										MUX_10_1_IN_4 => UNWINDOWED_692 ,
										MUX_10_1_IN_5 => UNWINDOWED_661 ,
										MUX_10_1_IN_6 => UNWINDOWED_724 ,
										MUX_10_1_IN_7 => UNWINDOWED_597 ,
										MUX_10_1_IN_8 => UNWINDOWED_852 ,
										MUX_10_1_IN_9 => UNWINDOWED_341 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_682
									);
MUX_REORD_UNIT_683 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_683 ,
										MUX_10_1_IN_1 => UNWINDOWED_683 ,
										MUX_10_1_IN_2 => UNWINDOWED_686 ,
										MUX_10_1_IN_3 => UNWINDOWED_679 ,
										MUX_10_1_IN_4 => UNWINDOWED_694 ,
										MUX_10_1_IN_5 => UNWINDOWED_663 ,
										MUX_10_1_IN_6 => UNWINDOWED_726 ,
										MUX_10_1_IN_7 => UNWINDOWED_599 ,
										MUX_10_1_IN_8 => UNWINDOWED_854 ,
										MUX_10_1_IN_9 => UNWINDOWED_343 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_683
									);
MUX_REORD_UNIT_684 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_684 ,
										MUX_10_1_IN_1 => UNWINDOWED_684 ,
										MUX_10_1_IN_2 => UNWINDOWED_681 ,
										MUX_10_1_IN_3 => UNWINDOWED_681 ,
										MUX_10_1_IN_4 => UNWINDOWED_696 ,
										MUX_10_1_IN_5 => UNWINDOWED_665 ,
										MUX_10_1_IN_6 => UNWINDOWED_728 ,
										MUX_10_1_IN_7 => UNWINDOWED_601 ,
										MUX_10_1_IN_8 => UNWINDOWED_856 ,
										MUX_10_1_IN_9 => UNWINDOWED_345 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_684
									);
MUX_REORD_UNIT_685 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_685 ,
										MUX_10_1_IN_1 => UNWINDOWED_686 ,
										MUX_10_1_IN_2 => UNWINDOWED_683 ,
										MUX_10_1_IN_3 => UNWINDOWED_683 ,
										MUX_10_1_IN_4 => UNWINDOWED_698 ,
										MUX_10_1_IN_5 => UNWINDOWED_667 ,
										MUX_10_1_IN_6 => UNWINDOWED_730 ,
										MUX_10_1_IN_7 => UNWINDOWED_603 ,
										MUX_10_1_IN_8 => UNWINDOWED_858 ,
										MUX_10_1_IN_9 => UNWINDOWED_347 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_685
									);
MUX_REORD_UNIT_686 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_686 ,
										MUX_10_1_IN_1 => UNWINDOWED_685 ,
										MUX_10_1_IN_2 => UNWINDOWED_685 ,
										MUX_10_1_IN_3 => UNWINDOWED_685 ,
										MUX_10_1_IN_4 => UNWINDOWED_700 ,
										MUX_10_1_IN_5 => UNWINDOWED_669 ,
										MUX_10_1_IN_6 => UNWINDOWED_732 ,
										MUX_10_1_IN_7 => UNWINDOWED_605 ,
										MUX_10_1_IN_8 => UNWINDOWED_860 ,
										MUX_10_1_IN_9 => UNWINDOWED_349 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_686
									);
MUX_REORD_UNIT_687 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_687 ,
										MUX_10_1_IN_1 => UNWINDOWED_687 ,
										MUX_10_1_IN_2 => UNWINDOWED_687 ,
										MUX_10_1_IN_3 => UNWINDOWED_687 ,
										MUX_10_1_IN_4 => UNWINDOWED_702 ,
										MUX_10_1_IN_5 => UNWINDOWED_671 ,
										MUX_10_1_IN_6 => UNWINDOWED_734 ,
										MUX_10_1_IN_7 => UNWINDOWED_607 ,
										MUX_10_1_IN_8 => UNWINDOWED_862 ,
										MUX_10_1_IN_9 => UNWINDOWED_351 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_687
									);
MUX_REORD_UNIT_688 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_688 ,
										MUX_10_1_IN_1 => UNWINDOWED_688 ,
										MUX_10_1_IN_2 => UNWINDOWED_688 ,
										MUX_10_1_IN_3 => UNWINDOWED_688 ,
										MUX_10_1_IN_4 => UNWINDOWED_673 ,
										MUX_10_1_IN_5 => UNWINDOWED_673 ,
										MUX_10_1_IN_6 => UNWINDOWED_736 ,
										MUX_10_1_IN_7 => UNWINDOWED_609 ,
										MUX_10_1_IN_8 => UNWINDOWED_864 ,
										MUX_10_1_IN_9 => UNWINDOWED_353 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_688
									);
MUX_REORD_UNIT_689 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_689 ,
										MUX_10_1_IN_1 => UNWINDOWED_690 ,
										MUX_10_1_IN_2 => UNWINDOWED_690 ,
										MUX_10_1_IN_3 => UNWINDOWED_690 ,
										MUX_10_1_IN_4 => UNWINDOWED_675 ,
										MUX_10_1_IN_5 => UNWINDOWED_675 ,
										MUX_10_1_IN_6 => UNWINDOWED_738 ,
										MUX_10_1_IN_7 => UNWINDOWED_611 ,
										MUX_10_1_IN_8 => UNWINDOWED_866 ,
										MUX_10_1_IN_9 => UNWINDOWED_355 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_689
									);
MUX_REORD_UNIT_690 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_690 ,
										MUX_10_1_IN_1 => UNWINDOWED_689 ,
										MUX_10_1_IN_2 => UNWINDOWED_692 ,
										MUX_10_1_IN_3 => UNWINDOWED_692 ,
										MUX_10_1_IN_4 => UNWINDOWED_677 ,
										MUX_10_1_IN_5 => UNWINDOWED_677 ,
										MUX_10_1_IN_6 => UNWINDOWED_740 ,
										MUX_10_1_IN_7 => UNWINDOWED_613 ,
										MUX_10_1_IN_8 => UNWINDOWED_868 ,
										MUX_10_1_IN_9 => UNWINDOWED_357 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_690
									);
MUX_REORD_UNIT_691 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_691 ,
										MUX_10_1_IN_1 => UNWINDOWED_691 ,
										MUX_10_1_IN_2 => UNWINDOWED_694 ,
										MUX_10_1_IN_3 => UNWINDOWED_694 ,
										MUX_10_1_IN_4 => UNWINDOWED_679 ,
										MUX_10_1_IN_5 => UNWINDOWED_679 ,
										MUX_10_1_IN_6 => UNWINDOWED_742 ,
										MUX_10_1_IN_7 => UNWINDOWED_615 ,
										MUX_10_1_IN_8 => UNWINDOWED_870 ,
										MUX_10_1_IN_9 => UNWINDOWED_359 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_691
									);
MUX_REORD_UNIT_692 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_692 ,
										MUX_10_1_IN_1 => UNWINDOWED_692 ,
										MUX_10_1_IN_2 => UNWINDOWED_689 ,
										MUX_10_1_IN_3 => UNWINDOWED_696 ,
										MUX_10_1_IN_4 => UNWINDOWED_681 ,
										MUX_10_1_IN_5 => UNWINDOWED_681 ,
										MUX_10_1_IN_6 => UNWINDOWED_744 ,
										MUX_10_1_IN_7 => UNWINDOWED_617 ,
										MUX_10_1_IN_8 => UNWINDOWED_872 ,
										MUX_10_1_IN_9 => UNWINDOWED_361 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_692
									);
MUX_REORD_UNIT_693 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_693 ,
										MUX_10_1_IN_1 => UNWINDOWED_694 ,
										MUX_10_1_IN_2 => UNWINDOWED_691 ,
										MUX_10_1_IN_3 => UNWINDOWED_698 ,
										MUX_10_1_IN_4 => UNWINDOWED_683 ,
										MUX_10_1_IN_5 => UNWINDOWED_683 ,
										MUX_10_1_IN_6 => UNWINDOWED_746 ,
										MUX_10_1_IN_7 => UNWINDOWED_619 ,
										MUX_10_1_IN_8 => UNWINDOWED_874 ,
										MUX_10_1_IN_9 => UNWINDOWED_363 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_693
									);
MUX_REORD_UNIT_694 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_694 ,
										MUX_10_1_IN_1 => UNWINDOWED_693 ,
										MUX_10_1_IN_2 => UNWINDOWED_693 ,
										MUX_10_1_IN_3 => UNWINDOWED_700 ,
										MUX_10_1_IN_4 => UNWINDOWED_685 ,
										MUX_10_1_IN_5 => UNWINDOWED_685 ,
										MUX_10_1_IN_6 => UNWINDOWED_748 ,
										MUX_10_1_IN_7 => UNWINDOWED_621 ,
										MUX_10_1_IN_8 => UNWINDOWED_876 ,
										MUX_10_1_IN_9 => UNWINDOWED_365 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_694
									);
MUX_REORD_UNIT_695 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_695 ,
										MUX_10_1_IN_1 => UNWINDOWED_695 ,
										MUX_10_1_IN_2 => UNWINDOWED_695 ,
										MUX_10_1_IN_3 => UNWINDOWED_702 ,
										MUX_10_1_IN_4 => UNWINDOWED_687 ,
										MUX_10_1_IN_5 => UNWINDOWED_687 ,
										MUX_10_1_IN_6 => UNWINDOWED_750 ,
										MUX_10_1_IN_7 => UNWINDOWED_623 ,
										MUX_10_1_IN_8 => UNWINDOWED_878 ,
										MUX_10_1_IN_9 => UNWINDOWED_367 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_695
									);
MUX_REORD_UNIT_696 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_696 ,
										MUX_10_1_IN_1 => UNWINDOWED_696 ,
										MUX_10_1_IN_2 => UNWINDOWED_696 ,
										MUX_10_1_IN_3 => UNWINDOWED_689 ,
										MUX_10_1_IN_4 => UNWINDOWED_689 ,
										MUX_10_1_IN_5 => UNWINDOWED_689 ,
										MUX_10_1_IN_6 => UNWINDOWED_752 ,
										MUX_10_1_IN_7 => UNWINDOWED_625 ,
										MUX_10_1_IN_8 => UNWINDOWED_880 ,
										MUX_10_1_IN_9 => UNWINDOWED_369 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_696
									);
MUX_REORD_UNIT_697 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_697 ,
										MUX_10_1_IN_1 => UNWINDOWED_698 ,
										MUX_10_1_IN_2 => UNWINDOWED_698 ,
										MUX_10_1_IN_3 => UNWINDOWED_691 ,
										MUX_10_1_IN_4 => UNWINDOWED_691 ,
										MUX_10_1_IN_5 => UNWINDOWED_691 ,
										MUX_10_1_IN_6 => UNWINDOWED_754 ,
										MUX_10_1_IN_7 => UNWINDOWED_627 ,
										MUX_10_1_IN_8 => UNWINDOWED_882 ,
										MUX_10_1_IN_9 => UNWINDOWED_371 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_697
									);
MUX_REORD_UNIT_698 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_698 ,
										MUX_10_1_IN_1 => UNWINDOWED_697 ,
										MUX_10_1_IN_2 => UNWINDOWED_700 ,
										MUX_10_1_IN_3 => UNWINDOWED_693 ,
										MUX_10_1_IN_4 => UNWINDOWED_693 ,
										MUX_10_1_IN_5 => UNWINDOWED_693 ,
										MUX_10_1_IN_6 => UNWINDOWED_756 ,
										MUX_10_1_IN_7 => UNWINDOWED_629 ,
										MUX_10_1_IN_8 => UNWINDOWED_884 ,
										MUX_10_1_IN_9 => UNWINDOWED_373 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_698
									);
MUX_REORD_UNIT_699 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_699 ,
										MUX_10_1_IN_1 => UNWINDOWED_699 ,
										MUX_10_1_IN_2 => UNWINDOWED_702 ,
										MUX_10_1_IN_3 => UNWINDOWED_695 ,
										MUX_10_1_IN_4 => UNWINDOWED_695 ,
										MUX_10_1_IN_5 => UNWINDOWED_695 ,
										MUX_10_1_IN_6 => UNWINDOWED_758 ,
										MUX_10_1_IN_7 => UNWINDOWED_631 ,
										MUX_10_1_IN_8 => UNWINDOWED_886 ,
										MUX_10_1_IN_9 => UNWINDOWED_375 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_699
									);
MUX_REORD_UNIT_700 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_700 ,
										MUX_10_1_IN_1 => UNWINDOWED_700 ,
										MUX_10_1_IN_2 => UNWINDOWED_697 ,
										MUX_10_1_IN_3 => UNWINDOWED_697 ,
										MUX_10_1_IN_4 => UNWINDOWED_697 ,
										MUX_10_1_IN_5 => UNWINDOWED_697 ,
										MUX_10_1_IN_6 => UNWINDOWED_760 ,
										MUX_10_1_IN_7 => UNWINDOWED_633 ,
										MUX_10_1_IN_8 => UNWINDOWED_888 ,
										MUX_10_1_IN_9 => UNWINDOWED_377 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_700
									);
MUX_REORD_UNIT_701 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_701 ,
										MUX_10_1_IN_1 => UNWINDOWED_702 ,
										MUX_10_1_IN_2 => UNWINDOWED_699 ,
										MUX_10_1_IN_3 => UNWINDOWED_699 ,
										MUX_10_1_IN_4 => UNWINDOWED_699 ,
										MUX_10_1_IN_5 => UNWINDOWED_699 ,
										MUX_10_1_IN_6 => UNWINDOWED_762 ,
										MUX_10_1_IN_7 => UNWINDOWED_635 ,
										MUX_10_1_IN_8 => UNWINDOWED_890 ,
										MUX_10_1_IN_9 => UNWINDOWED_379 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_701
									);
MUX_REORD_UNIT_702 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_702 ,
										MUX_10_1_IN_1 => UNWINDOWED_701 ,
										MUX_10_1_IN_2 => UNWINDOWED_701 ,
										MUX_10_1_IN_3 => UNWINDOWED_701 ,
										MUX_10_1_IN_4 => UNWINDOWED_701 ,
										MUX_10_1_IN_5 => UNWINDOWED_701 ,
										MUX_10_1_IN_6 => UNWINDOWED_764 ,
										MUX_10_1_IN_7 => UNWINDOWED_637 ,
										MUX_10_1_IN_8 => UNWINDOWED_892 ,
										MUX_10_1_IN_9 => UNWINDOWED_381 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_702
									);
MUX_REORD_UNIT_703 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_703 ,
										MUX_10_1_IN_1 => UNWINDOWED_703 ,
										MUX_10_1_IN_2 => UNWINDOWED_703 ,
										MUX_10_1_IN_3 => UNWINDOWED_703 ,
										MUX_10_1_IN_4 => UNWINDOWED_703 ,
										MUX_10_1_IN_5 => UNWINDOWED_703 ,
										MUX_10_1_IN_6 => UNWINDOWED_766 ,
										MUX_10_1_IN_7 => UNWINDOWED_639 ,
										MUX_10_1_IN_8 => UNWINDOWED_894 ,
										MUX_10_1_IN_9 => UNWINDOWED_383 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_703
									);
MUX_REORD_UNIT_704 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_704 ,
										MUX_10_1_IN_1 => UNWINDOWED_704 ,
										MUX_10_1_IN_2 => UNWINDOWED_704 ,
										MUX_10_1_IN_3 => UNWINDOWED_704 ,
										MUX_10_1_IN_4 => UNWINDOWED_704 ,
										MUX_10_1_IN_5 => UNWINDOWED_704 ,
										MUX_10_1_IN_6 => UNWINDOWED_641 ,
										MUX_10_1_IN_7 => UNWINDOWED_641 ,
										MUX_10_1_IN_8 => UNWINDOWED_896 ,
										MUX_10_1_IN_9 => UNWINDOWED_385 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_704
									);
MUX_REORD_UNIT_705 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_705 ,
										MUX_10_1_IN_1 => UNWINDOWED_706 ,
										MUX_10_1_IN_2 => UNWINDOWED_706 ,
										MUX_10_1_IN_3 => UNWINDOWED_706 ,
										MUX_10_1_IN_4 => UNWINDOWED_706 ,
										MUX_10_1_IN_5 => UNWINDOWED_706 ,
										MUX_10_1_IN_6 => UNWINDOWED_643 ,
										MUX_10_1_IN_7 => UNWINDOWED_643 ,
										MUX_10_1_IN_8 => UNWINDOWED_898 ,
										MUX_10_1_IN_9 => UNWINDOWED_387 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_705
									);
MUX_REORD_UNIT_706 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_706 ,
										MUX_10_1_IN_1 => UNWINDOWED_705 ,
										MUX_10_1_IN_2 => UNWINDOWED_708 ,
										MUX_10_1_IN_3 => UNWINDOWED_708 ,
										MUX_10_1_IN_4 => UNWINDOWED_708 ,
										MUX_10_1_IN_5 => UNWINDOWED_708 ,
										MUX_10_1_IN_6 => UNWINDOWED_645 ,
										MUX_10_1_IN_7 => UNWINDOWED_645 ,
										MUX_10_1_IN_8 => UNWINDOWED_900 ,
										MUX_10_1_IN_9 => UNWINDOWED_389 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_706
									);
MUX_REORD_UNIT_707 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_707 ,
										MUX_10_1_IN_1 => UNWINDOWED_707 ,
										MUX_10_1_IN_2 => UNWINDOWED_710 ,
										MUX_10_1_IN_3 => UNWINDOWED_710 ,
										MUX_10_1_IN_4 => UNWINDOWED_710 ,
										MUX_10_1_IN_5 => UNWINDOWED_710 ,
										MUX_10_1_IN_6 => UNWINDOWED_647 ,
										MUX_10_1_IN_7 => UNWINDOWED_647 ,
										MUX_10_1_IN_8 => UNWINDOWED_902 ,
										MUX_10_1_IN_9 => UNWINDOWED_391 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_707
									);
MUX_REORD_UNIT_708 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_708 ,
										MUX_10_1_IN_1 => UNWINDOWED_708 ,
										MUX_10_1_IN_2 => UNWINDOWED_705 ,
										MUX_10_1_IN_3 => UNWINDOWED_712 ,
										MUX_10_1_IN_4 => UNWINDOWED_712 ,
										MUX_10_1_IN_5 => UNWINDOWED_712 ,
										MUX_10_1_IN_6 => UNWINDOWED_649 ,
										MUX_10_1_IN_7 => UNWINDOWED_649 ,
										MUX_10_1_IN_8 => UNWINDOWED_904 ,
										MUX_10_1_IN_9 => UNWINDOWED_393 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_708
									);
MUX_REORD_UNIT_709 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_709 ,
										MUX_10_1_IN_1 => UNWINDOWED_710 ,
										MUX_10_1_IN_2 => UNWINDOWED_707 ,
										MUX_10_1_IN_3 => UNWINDOWED_714 ,
										MUX_10_1_IN_4 => UNWINDOWED_714 ,
										MUX_10_1_IN_5 => UNWINDOWED_714 ,
										MUX_10_1_IN_6 => UNWINDOWED_651 ,
										MUX_10_1_IN_7 => UNWINDOWED_651 ,
										MUX_10_1_IN_8 => UNWINDOWED_906 ,
										MUX_10_1_IN_9 => UNWINDOWED_395 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_709
									);
MUX_REORD_UNIT_710 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_710 ,
										MUX_10_1_IN_1 => UNWINDOWED_709 ,
										MUX_10_1_IN_2 => UNWINDOWED_709 ,
										MUX_10_1_IN_3 => UNWINDOWED_716 ,
										MUX_10_1_IN_4 => UNWINDOWED_716 ,
										MUX_10_1_IN_5 => UNWINDOWED_716 ,
										MUX_10_1_IN_6 => UNWINDOWED_653 ,
										MUX_10_1_IN_7 => UNWINDOWED_653 ,
										MUX_10_1_IN_8 => UNWINDOWED_908 ,
										MUX_10_1_IN_9 => UNWINDOWED_397 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_710
									);
MUX_REORD_UNIT_711 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_711 ,
										MUX_10_1_IN_1 => UNWINDOWED_711 ,
										MUX_10_1_IN_2 => UNWINDOWED_711 ,
										MUX_10_1_IN_3 => UNWINDOWED_718 ,
										MUX_10_1_IN_4 => UNWINDOWED_718 ,
										MUX_10_1_IN_5 => UNWINDOWED_718 ,
										MUX_10_1_IN_6 => UNWINDOWED_655 ,
										MUX_10_1_IN_7 => UNWINDOWED_655 ,
										MUX_10_1_IN_8 => UNWINDOWED_910 ,
										MUX_10_1_IN_9 => UNWINDOWED_399 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_711
									);
MUX_REORD_UNIT_712 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_712 ,
										MUX_10_1_IN_1 => UNWINDOWED_712 ,
										MUX_10_1_IN_2 => UNWINDOWED_712 ,
										MUX_10_1_IN_3 => UNWINDOWED_705 ,
										MUX_10_1_IN_4 => UNWINDOWED_720 ,
										MUX_10_1_IN_5 => UNWINDOWED_720 ,
										MUX_10_1_IN_6 => UNWINDOWED_657 ,
										MUX_10_1_IN_7 => UNWINDOWED_657 ,
										MUX_10_1_IN_8 => UNWINDOWED_912 ,
										MUX_10_1_IN_9 => UNWINDOWED_401 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_712
									);
MUX_REORD_UNIT_713 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_713 ,
										MUX_10_1_IN_1 => UNWINDOWED_714 ,
										MUX_10_1_IN_2 => UNWINDOWED_714 ,
										MUX_10_1_IN_3 => UNWINDOWED_707 ,
										MUX_10_1_IN_4 => UNWINDOWED_722 ,
										MUX_10_1_IN_5 => UNWINDOWED_722 ,
										MUX_10_1_IN_6 => UNWINDOWED_659 ,
										MUX_10_1_IN_7 => UNWINDOWED_659 ,
										MUX_10_1_IN_8 => UNWINDOWED_914 ,
										MUX_10_1_IN_9 => UNWINDOWED_403 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_713
									);
MUX_REORD_UNIT_714 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_714 ,
										MUX_10_1_IN_1 => UNWINDOWED_713 ,
										MUX_10_1_IN_2 => UNWINDOWED_716 ,
										MUX_10_1_IN_3 => UNWINDOWED_709 ,
										MUX_10_1_IN_4 => UNWINDOWED_724 ,
										MUX_10_1_IN_5 => UNWINDOWED_724 ,
										MUX_10_1_IN_6 => UNWINDOWED_661 ,
										MUX_10_1_IN_7 => UNWINDOWED_661 ,
										MUX_10_1_IN_8 => UNWINDOWED_916 ,
										MUX_10_1_IN_9 => UNWINDOWED_405 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_714
									);
MUX_REORD_UNIT_715 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_715 ,
										MUX_10_1_IN_1 => UNWINDOWED_715 ,
										MUX_10_1_IN_2 => UNWINDOWED_718 ,
										MUX_10_1_IN_3 => UNWINDOWED_711 ,
										MUX_10_1_IN_4 => UNWINDOWED_726 ,
										MUX_10_1_IN_5 => UNWINDOWED_726 ,
										MUX_10_1_IN_6 => UNWINDOWED_663 ,
										MUX_10_1_IN_7 => UNWINDOWED_663 ,
										MUX_10_1_IN_8 => UNWINDOWED_918 ,
										MUX_10_1_IN_9 => UNWINDOWED_407 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_715
									);
MUX_REORD_UNIT_716 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_716 ,
										MUX_10_1_IN_1 => UNWINDOWED_716 ,
										MUX_10_1_IN_2 => UNWINDOWED_713 ,
										MUX_10_1_IN_3 => UNWINDOWED_713 ,
										MUX_10_1_IN_4 => UNWINDOWED_728 ,
										MUX_10_1_IN_5 => UNWINDOWED_728 ,
										MUX_10_1_IN_6 => UNWINDOWED_665 ,
										MUX_10_1_IN_7 => UNWINDOWED_665 ,
										MUX_10_1_IN_8 => UNWINDOWED_920 ,
										MUX_10_1_IN_9 => UNWINDOWED_409 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_716
									);
MUX_REORD_UNIT_717 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_717 ,
										MUX_10_1_IN_1 => UNWINDOWED_718 ,
										MUX_10_1_IN_2 => UNWINDOWED_715 ,
										MUX_10_1_IN_3 => UNWINDOWED_715 ,
										MUX_10_1_IN_4 => UNWINDOWED_730 ,
										MUX_10_1_IN_5 => UNWINDOWED_730 ,
										MUX_10_1_IN_6 => UNWINDOWED_667 ,
										MUX_10_1_IN_7 => UNWINDOWED_667 ,
										MUX_10_1_IN_8 => UNWINDOWED_922 ,
										MUX_10_1_IN_9 => UNWINDOWED_411 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_717
									);
MUX_REORD_UNIT_718 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_718 ,
										MUX_10_1_IN_1 => UNWINDOWED_717 ,
										MUX_10_1_IN_2 => UNWINDOWED_717 ,
										MUX_10_1_IN_3 => UNWINDOWED_717 ,
										MUX_10_1_IN_4 => UNWINDOWED_732 ,
										MUX_10_1_IN_5 => UNWINDOWED_732 ,
										MUX_10_1_IN_6 => UNWINDOWED_669 ,
										MUX_10_1_IN_7 => UNWINDOWED_669 ,
										MUX_10_1_IN_8 => UNWINDOWED_924 ,
										MUX_10_1_IN_9 => UNWINDOWED_413 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_718
									);
MUX_REORD_UNIT_719 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_719 ,
										MUX_10_1_IN_1 => UNWINDOWED_719 ,
										MUX_10_1_IN_2 => UNWINDOWED_719 ,
										MUX_10_1_IN_3 => UNWINDOWED_719 ,
										MUX_10_1_IN_4 => UNWINDOWED_734 ,
										MUX_10_1_IN_5 => UNWINDOWED_734 ,
										MUX_10_1_IN_6 => UNWINDOWED_671 ,
										MUX_10_1_IN_7 => UNWINDOWED_671 ,
										MUX_10_1_IN_8 => UNWINDOWED_926 ,
										MUX_10_1_IN_9 => UNWINDOWED_415 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_719
									);
MUX_REORD_UNIT_720 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_720 ,
										MUX_10_1_IN_1 => UNWINDOWED_720 ,
										MUX_10_1_IN_2 => UNWINDOWED_720 ,
										MUX_10_1_IN_3 => UNWINDOWED_720 ,
										MUX_10_1_IN_4 => UNWINDOWED_705 ,
										MUX_10_1_IN_5 => UNWINDOWED_736 ,
										MUX_10_1_IN_6 => UNWINDOWED_673 ,
										MUX_10_1_IN_7 => UNWINDOWED_673 ,
										MUX_10_1_IN_8 => UNWINDOWED_928 ,
										MUX_10_1_IN_9 => UNWINDOWED_417 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_720
									);
MUX_REORD_UNIT_721 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_721 ,
										MUX_10_1_IN_1 => UNWINDOWED_722 ,
										MUX_10_1_IN_2 => UNWINDOWED_722 ,
										MUX_10_1_IN_3 => UNWINDOWED_722 ,
										MUX_10_1_IN_4 => UNWINDOWED_707 ,
										MUX_10_1_IN_5 => UNWINDOWED_738 ,
										MUX_10_1_IN_6 => UNWINDOWED_675 ,
										MUX_10_1_IN_7 => UNWINDOWED_675 ,
										MUX_10_1_IN_8 => UNWINDOWED_930 ,
										MUX_10_1_IN_9 => UNWINDOWED_419 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_721
									);
MUX_REORD_UNIT_722 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_722 ,
										MUX_10_1_IN_1 => UNWINDOWED_721 ,
										MUX_10_1_IN_2 => UNWINDOWED_724 ,
										MUX_10_1_IN_3 => UNWINDOWED_724 ,
										MUX_10_1_IN_4 => UNWINDOWED_709 ,
										MUX_10_1_IN_5 => UNWINDOWED_740 ,
										MUX_10_1_IN_6 => UNWINDOWED_677 ,
										MUX_10_1_IN_7 => UNWINDOWED_677 ,
										MUX_10_1_IN_8 => UNWINDOWED_932 ,
										MUX_10_1_IN_9 => UNWINDOWED_421 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_722
									);
MUX_REORD_UNIT_723 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_723 ,
										MUX_10_1_IN_1 => UNWINDOWED_723 ,
										MUX_10_1_IN_2 => UNWINDOWED_726 ,
										MUX_10_1_IN_3 => UNWINDOWED_726 ,
										MUX_10_1_IN_4 => UNWINDOWED_711 ,
										MUX_10_1_IN_5 => UNWINDOWED_742 ,
										MUX_10_1_IN_6 => UNWINDOWED_679 ,
										MUX_10_1_IN_7 => UNWINDOWED_679 ,
										MUX_10_1_IN_8 => UNWINDOWED_934 ,
										MUX_10_1_IN_9 => UNWINDOWED_423 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_723
									);
MUX_REORD_UNIT_724 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_724 ,
										MUX_10_1_IN_1 => UNWINDOWED_724 ,
										MUX_10_1_IN_2 => UNWINDOWED_721 ,
										MUX_10_1_IN_3 => UNWINDOWED_728 ,
										MUX_10_1_IN_4 => UNWINDOWED_713 ,
										MUX_10_1_IN_5 => UNWINDOWED_744 ,
										MUX_10_1_IN_6 => UNWINDOWED_681 ,
										MUX_10_1_IN_7 => UNWINDOWED_681 ,
										MUX_10_1_IN_8 => UNWINDOWED_936 ,
										MUX_10_1_IN_9 => UNWINDOWED_425 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_724
									);
MUX_REORD_UNIT_725 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_725 ,
										MUX_10_1_IN_1 => UNWINDOWED_726 ,
										MUX_10_1_IN_2 => UNWINDOWED_723 ,
										MUX_10_1_IN_3 => UNWINDOWED_730 ,
										MUX_10_1_IN_4 => UNWINDOWED_715 ,
										MUX_10_1_IN_5 => UNWINDOWED_746 ,
										MUX_10_1_IN_6 => UNWINDOWED_683 ,
										MUX_10_1_IN_7 => UNWINDOWED_683 ,
										MUX_10_1_IN_8 => UNWINDOWED_938 ,
										MUX_10_1_IN_9 => UNWINDOWED_427 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_725
									);
MUX_REORD_UNIT_726 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_726 ,
										MUX_10_1_IN_1 => UNWINDOWED_725 ,
										MUX_10_1_IN_2 => UNWINDOWED_725 ,
										MUX_10_1_IN_3 => UNWINDOWED_732 ,
										MUX_10_1_IN_4 => UNWINDOWED_717 ,
										MUX_10_1_IN_5 => UNWINDOWED_748 ,
										MUX_10_1_IN_6 => UNWINDOWED_685 ,
										MUX_10_1_IN_7 => UNWINDOWED_685 ,
										MUX_10_1_IN_8 => UNWINDOWED_940 ,
										MUX_10_1_IN_9 => UNWINDOWED_429 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_726
									);
MUX_REORD_UNIT_727 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_727 ,
										MUX_10_1_IN_1 => UNWINDOWED_727 ,
										MUX_10_1_IN_2 => UNWINDOWED_727 ,
										MUX_10_1_IN_3 => UNWINDOWED_734 ,
										MUX_10_1_IN_4 => UNWINDOWED_719 ,
										MUX_10_1_IN_5 => UNWINDOWED_750 ,
										MUX_10_1_IN_6 => UNWINDOWED_687 ,
										MUX_10_1_IN_7 => UNWINDOWED_687 ,
										MUX_10_1_IN_8 => UNWINDOWED_942 ,
										MUX_10_1_IN_9 => UNWINDOWED_431 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_727
									);
MUX_REORD_UNIT_728 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_728 ,
										MUX_10_1_IN_1 => UNWINDOWED_728 ,
										MUX_10_1_IN_2 => UNWINDOWED_728 ,
										MUX_10_1_IN_3 => UNWINDOWED_721 ,
										MUX_10_1_IN_4 => UNWINDOWED_721 ,
										MUX_10_1_IN_5 => UNWINDOWED_752 ,
										MUX_10_1_IN_6 => UNWINDOWED_689 ,
										MUX_10_1_IN_7 => UNWINDOWED_689 ,
										MUX_10_1_IN_8 => UNWINDOWED_944 ,
										MUX_10_1_IN_9 => UNWINDOWED_433 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_728
									);
MUX_REORD_UNIT_729 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_729 ,
										MUX_10_1_IN_1 => UNWINDOWED_730 ,
										MUX_10_1_IN_2 => UNWINDOWED_730 ,
										MUX_10_1_IN_3 => UNWINDOWED_723 ,
										MUX_10_1_IN_4 => UNWINDOWED_723 ,
										MUX_10_1_IN_5 => UNWINDOWED_754 ,
										MUX_10_1_IN_6 => UNWINDOWED_691 ,
										MUX_10_1_IN_7 => UNWINDOWED_691 ,
										MUX_10_1_IN_8 => UNWINDOWED_946 ,
										MUX_10_1_IN_9 => UNWINDOWED_435 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_729
									);
MUX_REORD_UNIT_730 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_730 ,
										MUX_10_1_IN_1 => UNWINDOWED_729 ,
										MUX_10_1_IN_2 => UNWINDOWED_732 ,
										MUX_10_1_IN_3 => UNWINDOWED_725 ,
										MUX_10_1_IN_4 => UNWINDOWED_725 ,
										MUX_10_1_IN_5 => UNWINDOWED_756 ,
										MUX_10_1_IN_6 => UNWINDOWED_693 ,
										MUX_10_1_IN_7 => UNWINDOWED_693 ,
										MUX_10_1_IN_8 => UNWINDOWED_948 ,
										MUX_10_1_IN_9 => UNWINDOWED_437 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_730
									);
MUX_REORD_UNIT_731 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_731 ,
										MUX_10_1_IN_1 => UNWINDOWED_731 ,
										MUX_10_1_IN_2 => UNWINDOWED_734 ,
										MUX_10_1_IN_3 => UNWINDOWED_727 ,
										MUX_10_1_IN_4 => UNWINDOWED_727 ,
										MUX_10_1_IN_5 => UNWINDOWED_758 ,
										MUX_10_1_IN_6 => UNWINDOWED_695 ,
										MUX_10_1_IN_7 => UNWINDOWED_695 ,
										MUX_10_1_IN_8 => UNWINDOWED_950 ,
										MUX_10_1_IN_9 => UNWINDOWED_439 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_731
									);
MUX_REORD_UNIT_732 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_732 ,
										MUX_10_1_IN_1 => UNWINDOWED_732 ,
										MUX_10_1_IN_2 => UNWINDOWED_729 ,
										MUX_10_1_IN_3 => UNWINDOWED_729 ,
										MUX_10_1_IN_4 => UNWINDOWED_729 ,
										MUX_10_1_IN_5 => UNWINDOWED_760 ,
										MUX_10_1_IN_6 => UNWINDOWED_697 ,
										MUX_10_1_IN_7 => UNWINDOWED_697 ,
										MUX_10_1_IN_8 => UNWINDOWED_952 ,
										MUX_10_1_IN_9 => UNWINDOWED_441 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_732
									);
MUX_REORD_UNIT_733 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_733 ,
										MUX_10_1_IN_1 => UNWINDOWED_734 ,
										MUX_10_1_IN_2 => UNWINDOWED_731 ,
										MUX_10_1_IN_3 => UNWINDOWED_731 ,
										MUX_10_1_IN_4 => UNWINDOWED_731 ,
										MUX_10_1_IN_5 => UNWINDOWED_762 ,
										MUX_10_1_IN_6 => UNWINDOWED_699 ,
										MUX_10_1_IN_7 => UNWINDOWED_699 ,
										MUX_10_1_IN_8 => UNWINDOWED_954 ,
										MUX_10_1_IN_9 => UNWINDOWED_443 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_733
									);
MUX_REORD_UNIT_734 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_734 ,
										MUX_10_1_IN_1 => UNWINDOWED_733 ,
										MUX_10_1_IN_2 => UNWINDOWED_733 ,
										MUX_10_1_IN_3 => UNWINDOWED_733 ,
										MUX_10_1_IN_4 => UNWINDOWED_733 ,
										MUX_10_1_IN_5 => UNWINDOWED_764 ,
										MUX_10_1_IN_6 => UNWINDOWED_701 ,
										MUX_10_1_IN_7 => UNWINDOWED_701 ,
										MUX_10_1_IN_8 => UNWINDOWED_956 ,
										MUX_10_1_IN_9 => UNWINDOWED_445 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_734
									);
MUX_REORD_UNIT_735 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_735 ,
										MUX_10_1_IN_1 => UNWINDOWED_735 ,
										MUX_10_1_IN_2 => UNWINDOWED_735 ,
										MUX_10_1_IN_3 => UNWINDOWED_735 ,
										MUX_10_1_IN_4 => UNWINDOWED_735 ,
										MUX_10_1_IN_5 => UNWINDOWED_766 ,
										MUX_10_1_IN_6 => UNWINDOWED_703 ,
										MUX_10_1_IN_7 => UNWINDOWED_703 ,
										MUX_10_1_IN_8 => UNWINDOWED_958 ,
										MUX_10_1_IN_9 => UNWINDOWED_447 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_735
									);
MUX_REORD_UNIT_736 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_736 ,
										MUX_10_1_IN_1 => UNWINDOWED_736 ,
										MUX_10_1_IN_2 => UNWINDOWED_736 ,
										MUX_10_1_IN_3 => UNWINDOWED_736 ,
										MUX_10_1_IN_4 => UNWINDOWED_736 ,
										MUX_10_1_IN_5 => UNWINDOWED_705 ,
										MUX_10_1_IN_6 => UNWINDOWED_705 ,
										MUX_10_1_IN_7 => UNWINDOWED_705 ,
										MUX_10_1_IN_8 => UNWINDOWED_960 ,
										MUX_10_1_IN_9 => UNWINDOWED_449 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_736
									);
MUX_REORD_UNIT_737 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_737 ,
										MUX_10_1_IN_1 => UNWINDOWED_738 ,
										MUX_10_1_IN_2 => UNWINDOWED_738 ,
										MUX_10_1_IN_3 => UNWINDOWED_738 ,
										MUX_10_1_IN_4 => UNWINDOWED_738 ,
										MUX_10_1_IN_5 => UNWINDOWED_707 ,
										MUX_10_1_IN_6 => UNWINDOWED_707 ,
										MUX_10_1_IN_7 => UNWINDOWED_707 ,
										MUX_10_1_IN_8 => UNWINDOWED_962 ,
										MUX_10_1_IN_9 => UNWINDOWED_451 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_737
									);
MUX_REORD_UNIT_738 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_738 ,
										MUX_10_1_IN_1 => UNWINDOWED_737 ,
										MUX_10_1_IN_2 => UNWINDOWED_740 ,
										MUX_10_1_IN_3 => UNWINDOWED_740 ,
										MUX_10_1_IN_4 => UNWINDOWED_740 ,
										MUX_10_1_IN_5 => UNWINDOWED_709 ,
										MUX_10_1_IN_6 => UNWINDOWED_709 ,
										MUX_10_1_IN_7 => UNWINDOWED_709 ,
										MUX_10_1_IN_8 => UNWINDOWED_964 ,
										MUX_10_1_IN_9 => UNWINDOWED_453 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_738
									);
MUX_REORD_UNIT_739 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_739 ,
										MUX_10_1_IN_1 => UNWINDOWED_739 ,
										MUX_10_1_IN_2 => UNWINDOWED_742 ,
										MUX_10_1_IN_3 => UNWINDOWED_742 ,
										MUX_10_1_IN_4 => UNWINDOWED_742 ,
										MUX_10_1_IN_5 => UNWINDOWED_711 ,
										MUX_10_1_IN_6 => UNWINDOWED_711 ,
										MUX_10_1_IN_7 => UNWINDOWED_711 ,
										MUX_10_1_IN_8 => UNWINDOWED_966 ,
										MUX_10_1_IN_9 => UNWINDOWED_455 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_739
									);
MUX_REORD_UNIT_740 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_740 ,
										MUX_10_1_IN_1 => UNWINDOWED_740 ,
										MUX_10_1_IN_2 => UNWINDOWED_737 ,
										MUX_10_1_IN_3 => UNWINDOWED_744 ,
										MUX_10_1_IN_4 => UNWINDOWED_744 ,
										MUX_10_1_IN_5 => UNWINDOWED_713 ,
										MUX_10_1_IN_6 => UNWINDOWED_713 ,
										MUX_10_1_IN_7 => UNWINDOWED_713 ,
										MUX_10_1_IN_8 => UNWINDOWED_968 ,
										MUX_10_1_IN_9 => UNWINDOWED_457 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_740
									);
MUX_REORD_UNIT_741 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_741 ,
										MUX_10_1_IN_1 => UNWINDOWED_742 ,
										MUX_10_1_IN_2 => UNWINDOWED_739 ,
										MUX_10_1_IN_3 => UNWINDOWED_746 ,
										MUX_10_1_IN_4 => UNWINDOWED_746 ,
										MUX_10_1_IN_5 => UNWINDOWED_715 ,
										MUX_10_1_IN_6 => UNWINDOWED_715 ,
										MUX_10_1_IN_7 => UNWINDOWED_715 ,
										MUX_10_1_IN_8 => UNWINDOWED_970 ,
										MUX_10_1_IN_9 => UNWINDOWED_459 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_741
									);
MUX_REORD_UNIT_742 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_742 ,
										MUX_10_1_IN_1 => UNWINDOWED_741 ,
										MUX_10_1_IN_2 => UNWINDOWED_741 ,
										MUX_10_1_IN_3 => UNWINDOWED_748 ,
										MUX_10_1_IN_4 => UNWINDOWED_748 ,
										MUX_10_1_IN_5 => UNWINDOWED_717 ,
										MUX_10_1_IN_6 => UNWINDOWED_717 ,
										MUX_10_1_IN_7 => UNWINDOWED_717 ,
										MUX_10_1_IN_8 => UNWINDOWED_972 ,
										MUX_10_1_IN_9 => UNWINDOWED_461 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_742
									);
MUX_REORD_UNIT_743 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_743 ,
										MUX_10_1_IN_1 => UNWINDOWED_743 ,
										MUX_10_1_IN_2 => UNWINDOWED_743 ,
										MUX_10_1_IN_3 => UNWINDOWED_750 ,
										MUX_10_1_IN_4 => UNWINDOWED_750 ,
										MUX_10_1_IN_5 => UNWINDOWED_719 ,
										MUX_10_1_IN_6 => UNWINDOWED_719 ,
										MUX_10_1_IN_7 => UNWINDOWED_719 ,
										MUX_10_1_IN_8 => UNWINDOWED_974 ,
										MUX_10_1_IN_9 => UNWINDOWED_463 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_743
									);
MUX_REORD_UNIT_744 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_744 ,
										MUX_10_1_IN_1 => UNWINDOWED_744 ,
										MUX_10_1_IN_2 => UNWINDOWED_744 ,
										MUX_10_1_IN_3 => UNWINDOWED_737 ,
										MUX_10_1_IN_4 => UNWINDOWED_752 ,
										MUX_10_1_IN_5 => UNWINDOWED_721 ,
										MUX_10_1_IN_6 => UNWINDOWED_721 ,
										MUX_10_1_IN_7 => UNWINDOWED_721 ,
										MUX_10_1_IN_8 => UNWINDOWED_976 ,
										MUX_10_1_IN_9 => UNWINDOWED_465 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_744
									);
MUX_REORD_UNIT_745 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_745 ,
										MUX_10_1_IN_1 => UNWINDOWED_746 ,
										MUX_10_1_IN_2 => UNWINDOWED_746 ,
										MUX_10_1_IN_3 => UNWINDOWED_739 ,
										MUX_10_1_IN_4 => UNWINDOWED_754 ,
										MUX_10_1_IN_5 => UNWINDOWED_723 ,
										MUX_10_1_IN_6 => UNWINDOWED_723 ,
										MUX_10_1_IN_7 => UNWINDOWED_723 ,
										MUX_10_1_IN_8 => UNWINDOWED_978 ,
										MUX_10_1_IN_9 => UNWINDOWED_467 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_745
									);
MUX_REORD_UNIT_746 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_746 ,
										MUX_10_1_IN_1 => UNWINDOWED_745 ,
										MUX_10_1_IN_2 => UNWINDOWED_748 ,
										MUX_10_1_IN_3 => UNWINDOWED_741 ,
										MUX_10_1_IN_4 => UNWINDOWED_756 ,
										MUX_10_1_IN_5 => UNWINDOWED_725 ,
										MUX_10_1_IN_6 => UNWINDOWED_725 ,
										MUX_10_1_IN_7 => UNWINDOWED_725 ,
										MUX_10_1_IN_8 => UNWINDOWED_980 ,
										MUX_10_1_IN_9 => UNWINDOWED_469 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_746
									);
MUX_REORD_UNIT_747 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_747 ,
										MUX_10_1_IN_1 => UNWINDOWED_747 ,
										MUX_10_1_IN_2 => UNWINDOWED_750 ,
										MUX_10_1_IN_3 => UNWINDOWED_743 ,
										MUX_10_1_IN_4 => UNWINDOWED_758 ,
										MUX_10_1_IN_5 => UNWINDOWED_727 ,
										MUX_10_1_IN_6 => UNWINDOWED_727 ,
										MUX_10_1_IN_7 => UNWINDOWED_727 ,
										MUX_10_1_IN_8 => UNWINDOWED_982 ,
										MUX_10_1_IN_9 => UNWINDOWED_471 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_747
									);
MUX_REORD_UNIT_748 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_748 ,
										MUX_10_1_IN_1 => UNWINDOWED_748 ,
										MUX_10_1_IN_2 => UNWINDOWED_745 ,
										MUX_10_1_IN_3 => UNWINDOWED_745 ,
										MUX_10_1_IN_4 => UNWINDOWED_760 ,
										MUX_10_1_IN_5 => UNWINDOWED_729 ,
										MUX_10_1_IN_6 => UNWINDOWED_729 ,
										MUX_10_1_IN_7 => UNWINDOWED_729 ,
										MUX_10_1_IN_8 => UNWINDOWED_984 ,
										MUX_10_1_IN_9 => UNWINDOWED_473 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_748
									);
MUX_REORD_UNIT_749 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_749 ,
										MUX_10_1_IN_1 => UNWINDOWED_750 ,
										MUX_10_1_IN_2 => UNWINDOWED_747 ,
										MUX_10_1_IN_3 => UNWINDOWED_747 ,
										MUX_10_1_IN_4 => UNWINDOWED_762 ,
										MUX_10_1_IN_5 => UNWINDOWED_731 ,
										MUX_10_1_IN_6 => UNWINDOWED_731 ,
										MUX_10_1_IN_7 => UNWINDOWED_731 ,
										MUX_10_1_IN_8 => UNWINDOWED_986 ,
										MUX_10_1_IN_9 => UNWINDOWED_475 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_749
									);
MUX_REORD_UNIT_750 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_750 ,
										MUX_10_1_IN_1 => UNWINDOWED_749 ,
										MUX_10_1_IN_2 => UNWINDOWED_749 ,
										MUX_10_1_IN_3 => UNWINDOWED_749 ,
										MUX_10_1_IN_4 => UNWINDOWED_764 ,
										MUX_10_1_IN_5 => UNWINDOWED_733 ,
										MUX_10_1_IN_6 => UNWINDOWED_733 ,
										MUX_10_1_IN_7 => UNWINDOWED_733 ,
										MUX_10_1_IN_8 => UNWINDOWED_988 ,
										MUX_10_1_IN_9 => UNWINDOWED_477 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_750
									);
MUX_REORD_UNIT_751 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_751 ,
										MUX_10_1_IN_1 => UNWINDOWED_751 ,
										MUX_10_1_IN_2 => UNWINDOWED_751 ,
										MUX_10_1_IN_3 => UNWINDOWED_751 ,
										MUX_10_1_IN_4 => UNWINDOWED_766 ,
										MUX_10_1_IN_5 => UNWINDOWED_735 ,
										MUX_10_1_IN_6 => UNWINDOWED_735 ,
										MUX_10_1_IN_7 => UNWINDOWED_735 ,
										MUX_10_1_IN_8 => UNWINDOWED_990 ,
										MUX_10_1_IN_9 => UNWINDOWED_479 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_751
									);
MUX_REORD_UNIT_752 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_752 ,
										MUX_10_1_IN_1 => UNWINDOWED_752 ,
										MUX_10_1_IN_2 => UNWINDOWED_752 ,
										MUX_10_1_IN_3 => UNWINDOWED_752 ,
										MUX_10_1_IN_4 => UNWINDOWED_737 ,
										MUX_10_1_IN_5 => UNWINDOWED_737 ,
										MUX_10_1_IN_6 => UNWINDOWED_737 ,
										MUX_10_1_IN_7 => UNWINDOWED_737 ,
										MUX_10_1_IN_8 => UNWINDOWED_992 ,
										MUX_10_1_IN_9 => UNWINDOWED_481 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_752
									);
MUX_REORD_UNIT_753 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_753 ,
										MUX_10_1_IN_1 => UNWINDOWED_754 ,
										MUX_10_1_IN_2 => UNWINDOWED_754 ,
										MUX_10_1_IN_3 => UNWINDOWED_754 ,
										MUX_10_1_IN_4 => UNWINDOWED_739 ,
										MUX_10_1_IN_5 => UNWINDOWED_739 ,
										MUX_10_1_IN_6 => UNWINDOWED_739 ,
										MUX_10_1_IN_7 => UNWINDOWED_739 ,
										MUX_10_1_IN_8 => UNWINDOWED_994 ,
										MUX_10_1_IN_9 => UNWINDOWED_483 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_753
									);
MUX_REORD_UNIT_754 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_754 ,
										MUX_10_1_IN_1 => UNWINDOWED_753 ,
										MUX_10_1_IN_2 => UNWINDOWED_756 ,
										MUX_10_1_IN_3 => UNWINDOWED_756 ,
										MUX_10_1_IN_4 => UNWINDOWED_741 ,
										MUX_10_1_IN_5 => UNWINDOWED_741 ,
										MUX_10_1_IN_6 => UNWINDOWED_741 ,
										MUX_10_1_IN_7 => UNWINDOWED_741 ,
										MUX_10_1_IN_8 => UNWINDOWED_996 ,
										MUX_10_1_IN_9 => UNWINDOWED_485 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_754
									);
MUX_REORD_UNIT_755 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_755 ,
										MUX_10_1_IN_1 => UNWINDOWED_755 ,
										MUX_10_1_IN_2 => UNWINDOWED_758 ,
										MUX_10_1_IN_3 => UNWINDOWED_758 ,
										MUX_10_1_IN_4 => UNWINDOWED_743 ,
										MUX_10_1_IN_5 => UNWINDOWED_743 ,
										MUX_10_1_IN_6 => UNWINDOWED_743 ,
										MUX_10_1_IN_7 => UNWINDOWED_743 ,
										MUX_10_1_IN_8 => UNWINDOWED_998 ,
										MUX_10_1_IN_9 => UNWINDOWED_487 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_755
									);
MUX_REORD_UNIT_756 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_756 ,
										MUX_10_1_IN_1 => UNWINDOWED_756 ,
										MUX_10_1_IN_2 => UNWINDOWED_753 ,
										MUX_10_1_IN_3 => UNWINDOWED_760 ,
										MUX_10_1_IN_4 => UNWINDOWED_745 ,
										MUX_10_1_IN_5 => UNWINDOWED_745 ,
										MUX_10_1_IN_6 => UNWINDOWED_745 ,
										MUX_10_1_IN_7 => UNWINDOWED_745 ,
										MUX_10_1_IN_8 => UNWINDOWED_1000 ,
										MUX_10_1_IN_9 => UNWINDOWED_489 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_756
									);
MUX_REORD_UNIT_757 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_757 ,
										MUX_10_1_IN_1 => UNWINDOWED_758 ,
										MUX_10_1_IN_2 => UNWINDOWED_755 ,
										MUX_10_1_IN_3 => UNWINDOWED_762 ,
										MUX_10_1_IN_4 => UNWINDOWED_747 ,
										MUX_10_1_IN_5 => UNWINDOWED_747 ,
										MUX_10_1_IN_6 => UNWINDOWED_747 ,
										MUX_10_1_IN_7 => UNWINDOWED_747 ,
										MUX_10_1_IN_8 => UNWINDOWED_1002 ,
										MUX_10_1_IN_9 => UNWINDOWED_491 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_757
									);
MUX_REORD_UNIT_758 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_758 ,
										MUX_10_1_IN_1 => UNWINDOWED_757 ,
										MUX_10_1_IN_2 => UNWINDOWED_757 ,
										MUX_10_1_IN_3 => UNWINDOWED_764 ,
										MUX_10_1_IN_4 => UNWINDOWED_749 ,
										MUX_10_1_IN_5 => UNWINDOWED_749 ,
										MUX_10_1_IN_6 => UNWINDOWED_749 ,
										MUX_10_1_IN_7 => UNWINDOWED_749 ,
										MUX_10_1_IN_8 => UNWINDOWED_1004 ,
										MUX_10_1_IN_9 => UNWINDOWED_493 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_758
									);
MUX_REORD_UNIT_759 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_759 ,
										MUX_10_1_IN_1 => UNWINDOWED_759 ,
										MUX_10_1_IN_2 => UNWINDOWED_759 ,
										MUX_10_1_IN_3 => UNWINDOWED_766 ,
										MUX_10_1_IN_4 => UNWINDOWED_751 ,
										MUX_10_1_IN_5 => UNWINDOWED_751 ,
										MUX_10_1_IN_6 => UNWINDOWED_751 ,
										MUX_10_1_IN_7 => UNWINDOWED_751 ,
										MUX_10_1_IN_8 => UNWINDOWED_1006 ,
										MUX_10_1_IN_9 => UNWINDOWED_495 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_759
									);
MUX_REORD_UNIT_760 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_760 ,
										MUX_10_1_IN_1 => UNWINDOWED_760 ,
										MUX_10_1_IN_2 => UNWINDOWED_760 ,
										MUX_10_1_IN_3 => UNWINDOWED_753 ,
										MUX_10_1_IN_4 => UNWINDOWED_753 ,
										MUX_10_1_IN_5 => UNWINDOWED_753 ,
										MUX_10_1_IN_6 => UNWINDOWED_753 ,
										MUX_10_1_IN_7 => UNWINDOWED_753 ,
										MUX_10_1_IN_8 => UNWINDOWED_1008 ,
										MUX_10_1_IN_9 => UNWINDOWED_497 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_760
									);
MUX_REORD_UNIT_761 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_761 ,
										MUX_10_1_IN_1 => UNWINDOWED_762 ,
										MUX_10_1_IN_2 => UNWINDOWED_762 ,
										MUX_10_1_IN_3 => UNWINDOWED_755 ,
										MUX_10_1_IN_4 => UNWINDOWED_755 ,
										MUX_10_1_IN_5 => UNWINDOWED_755 ,
										MUX_10_1_IN_6 => UNWINDOWED_755 ,
										MUX_10_1_IN_7 => UNWINDOWED_755 ,
										MUX_10_1_IN_8 => UNWINDOWED_1010 ,
										MUX_10_1_IN_9 => UNWINDOWED_499 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_761
									);
MUX_REORD_UNIT_762 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_762 ,
										MUX_10_1_IN_1 => UNWINDOWED_761 ,
										MUX_10_1_IN_2 => UNWINDOWED_764 ,
										MUX_10_1_IN_3 => UNWINDOWED_757 ,
										MUX_10_1_IN_4 => UNWINDOWED_757 ,
										MUX_10_1_IN_5 => UNWINDOWED_757 ,
										MUX_10_1_IN_6 => UNWINDOWED_757 ,
										MUX_10_1_IN_7 => UNWINDOWED_757 ,
										MUX_10_1_IN_8 => UNWINDOWED_1012 ,
										MUX_10_1_IN_9 => UNWINDOWED_501 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_762
									);
MUX_REORD_UNIT_763 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_763 ,
										MUX_10_1_IN_1 => UNWINDOWED_763 ,
										MUX_10_1_IN_2 => UNWINDOWED_766 ,
										MUX_10_1_IN_3 => UNWINDOWED_759 ,
										MUX_10_1_IN_4 => UNWINDOWED_759 ,
										MUX_10_1_IN_5 => UNWINDOWED_759 ,
										MUX_10_1_IN_6 => UNWINDOWED_759 ,
										MUX_10_1_IN_7 => UNWINDOWED_759 ,
										MUX_10_1_IN_8 => UNWINDOWED_1014 ,
										MUX_10_1_IN_9 => UNWINDOWED_503 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_763
									);
MUX_REORD_UNIT_764 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_764 ,
										MUX_10_1_IN_1 => UNWINDOWED_764 ,
										MUX_10_1_IN_2 => UNWINDOWED_761 ,
										MUX_10_1_IN_3 => UNWINDOWED_761 ,
										MUX_10_1_IN_4 => UNWINDOWED_761 ,
										MUX_10_1_IN_5 => UNWINDOWED_761 ,
										MUX_10_1_IN_6 => UNWINDOWED_761 ,
										MUX_10_1_IN_7 => UNWINDOWED_761 ,
										MUX_10_1_IN_8 => UNWINDOWED_1016 ,
										MUX_10_1_IN_9 => UNWINDOWED_505 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_764
									);
MUX_REORD_UNIT_765 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_765 ,
										MUX_10_1_IN_1 => UNWINDOWED_766 ,
										MUX_10_1_IN_2 => UNWINDOWED_763 ,
										MUX_10_1_IN_3 => UNWINDOWED_763 ,
										MUX_10_1_IN_4 => UNWINDOWED_763 ,
										MUX_10_1_IN_5 => UNWINDOWED_763 ,
										MUX_10_1_IN_6 => UNWINDOWED_763 ,
										MUX_10_1_IN_7 => UNWINDOWED_763 ,
										MUX_10_1_IN_8 => UNWINDOWED_1018 ,
										MUX_10_1_IN_9 => UNWINDOWED_507 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_765
									);
MUX_REORD_UNIT_766 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_766 ,
										MUX_10_1_IN_1 => UNWINDOWED_765 ,
										MUX_10_1_IN_2 => UNWINDOWED_765 ,
										MUX_10_1_IN_3 => UNWINDOWED_765 ,
										MUX_10_1_IN_4 => UNWINDOWED_765 ,
										MUX_10_1_IN_5 => UNWINDOWED_765 ,
										MUX_10_1_IN_6 => UNWINDOWED_765 ,
										MUX_10_1_IN_7 => UNWINDOWED_765 ,
										MUX_10_1_IN_8 => UNWINDOWED_1020 ,
										MUX_10_1_IN_9 => UNWINDOWED_509 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_766
									);
MUX_REORD_UNIT_767 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_767 ,
										MUX_10_1_IN_1 => UNWINDOWED_767 ,
										MUX_10_1_IN_2 => UNWINDOWED_767 ,
										MUX_10_1_IN_3 => UNWINDOWED_767 ,
										MUX_10_1_IN_4 => UNWINDOWED_767 ,
										MUX_10_1_IN_5 => UNWINDOWED_767 ,
										MUX_10_1_IN_6 => UNWINDOWED_767 ,
										MUX_10_1_IN_7 => UNWINDOWED_767 ,
										MUX_10_1_IN_8 => UNWINDOWED_1022 ,
										MUX_10_1_IN_9 => UNWINDOWED_511 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_767
									);
MUX_REORD_UNIT_768 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_768 ,
										MUX_10_1_IN_1 => UNWINDOWED_768 ,
										MUX_10_1_IN_2 => UNWINDOWED_768 ,
										MUX_10_1_IN_3 => UNWINDOWED_768 ,
										MUX_10_1_IN_4 => UNWINDOWED_768 ,
										MUX_10_1_IN_5 => UNWINDOWED_768 ,
										MUX_10_1_IN_6 => UNWINDOWED_768 ,
										MUX_10_1_IN_7 => UNWINDOWED_768 ,
										MUX_10_1_IN_8 => UNWINDOWED_513 ,
										MUX_10_1_IN_9 => UNWINDOWED_513 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_768
									);
MUX_REORD_UNIT_769 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_769 ,
										MUX_10_1_IN_1 => UNWINDOWED_770 ,
										MUX_10_1_IN_2 => UNWINDOWED_770 ,
										MUX_10_1_IN_3 => UNWINDOWED_770 ,
										MUX_10_1_IN_4 => UNWINDOWED_770 ,
										MUX_10_1_IN_5 => UNWINDOWED_770 ,
										MUX_10_1_IN_6 => UNWINDOWED_770 ,
										MUX_10_1_IN_7 => UNWINDOWED_770 ,
										MUX_10_1_IN_8 => UNWINDOWED_515 ,
										MUX_10_1_IN_9 => UNWINDOWED_515 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_769
									);
MUX_REORD_UNIT_770 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_770 ,
										MUX_10_1_IN_1 => UNWINDOWED_769 ,
										MUX_10_1_IN_2 => UNWINDOWED_772 ,
										MUX_10_1_IN_3 => UNWINDOWED_772 ,
										MUX_10_1_IN_4 => UNWINDOWED_772 ,
										MUX_10_1_IN_5 => UNWINDOWED_772 ,
										MUX_10_1_IN_6 => UNWINDOWED_772 ,
										MUX_10_1_IN_7 => UNWINDOWED_772 ,
										MUX_10_1_IN_8 => UNWINDOWED_517 ,
										MUX_10_1_IN_9 => UNWINDOWED_517 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_770
									);
MUX_REORD_UNIT_771 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_771 ,
										MUX_10_1_IN_1 => UNWINDOWED_771 ,
										MUX_10_1_IN_2 => UNWINDOWED_774 ,
										MUX_10_1_IN_3 => UNWINDOWED_774 ,
										MUX_10_1_IN_4 => UNWINDOWED_774 ,
										MUX_10_1_IN_5 => UNWINDOWED_774 ,
										MUX_10_1_IN_6 => UNWINDOWED_774 ,
										MUX_10_1_IN_7 => UNWINDOWED_774 ,
										MUX_10_1_IN_8 => UNWINDOWED_519 ,
										MUX_10_1_IN_9 => UNWINDOWED_519 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_771
									);
MUX_REORD_UNIT_772 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_772 ,
										MUX_10_1_IN_1 => UNWINDOWED_772 ,
										MUX_10_1_IN_2 => UNWINDOWED_769 ,
										MUX_10_1_IN_3 => UNWINDOWED_776 ,
										MUX_10_1_IN_4 => UNWINDOWED_776 ,
										MUX_10_1_IN_5 => UNWINDOWED_776 ,
										MUX_10_1_IN_6 => UNWINDOWED_776 ,
										MUX_10_1_IN_7 => UNWINDOWED_776 ,
										MUX_10_1_IN_8 => UNWINDOWED_521 ,
										MUX_10_1_IN_9 => UNWINDOWED_521 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_772
									);
MUX_REORD_UNIT_773 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_773 ,
										MUX_10_1_IN_1 => UNWINDOWED_774 ,
										MUX_10_1_IN_2 => UNWINDOWED_771 ,
										MUX_10_1_IN_3 => UNWINDOWED_778 ,
										MUX_10_1_IN_4 => UNWINDOWED_778 ,
										MUX_10_1_IN_5 => UNWINDOWED_778 ,
										MUX_10_1_IN_6 => UNWINDOWED_778 ,
										MUX_10_1_IN_7 => UNWINDOWED_778 ,
										MUX_10_1_IN_8 => UNWINDOWED_523 ,
										MUX_10_1_IN_9 => UNWINDOWED_523 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_773
									);
MUX_REORD_UNIT_774 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_774 ,
										MUX_10_1_IN_1 => UNWINDOWED_773 ,
										MUX_10_1_IN_2 => UNWINDOWED_773 ,
										MUX_10_1_IN_3 => UNWINDOWED_780 ,
										MUX_10_1_IN_4 => UNWINDOWED_780 ,
										MUX_10_1_IN_5 => UNWINDOWED_780 ,
										MUX_10_1_IN_6 => UNWINDOWED_780 ,
										MUX_10_1_IN_7 => UNWINDOWED_780 ,
										MUX_10_1_IN_8 => UNWINDOWED_525 ,
										MUX_10_1_IN_9 => UNWINDOWED_525 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_774
									);
MUX_REORD_UNIT_775 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_775 ,
										MUX_10_1_IN_1 => UNWINDOWED_775 ,
										MUX_10_1_IN_2 => UNWINDOWED_775 ,
										MUX_10_1_IN_3 => UNWINDOWED_782 ,
										MUX_10_1_IN_4 => UNWINDOWED_782 ,
										MUX_10_1_IN_5 => UNWINDOWED_782 ,
										MUX_10_1_IN_6 => UNWINDOWED_782 ,
										MUX_10_1_IN_7 => UNWINDOWED_782 ,
										MUX_10_1_IN_8 => UNWINDOWED_527 ,
										MUX_10_1_IN_9 => UNWINDOWED_527 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_775
									);
MUX_REORD_UNIT_776 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_776 ,
										MUX_10_1_IN_1 => UNWINDOWED_776 ,
										MUX_10_1_IN_2 => UNWINDOWED_776 ,
										MUX_10_1_IN_3 => UNWINDOWED_769 ,
										MUX_10_1_IN_4 => UNWINDOWED_784 ,
										MUX_10_1_IN_5 => UNWINDOWED_784 ,
										MUX_10_1_IN_6 => UNWINDOWED_784 ,
										MUX_10_1_IN_7 => UNWINDOWED_784 ,
										MUX_10_1_IN_8 => UNWINDOWED_529 ,
										MUX_10_1_IN_9 => UNWINDOWED_529 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_776
									);
MUX_REORD_UNIT_777 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_777 ,
										MUX_10_1_IN_1 => UNWINDOWED_778 ,
										MUX_10_1_IN_2 => UNWINDOWED_778 ,
										MUX_10_1_IN_3 => UNWINDOWED_771 ,
										MUX_10_1_IN_4 => UNWINDOWED_786 ,
										MUX_10_1_IN_5 => UNWINDOWED_786 ,
										MUX_10_1_IN_6 => UNWINDOWED_786 ,
										MUX_10_1_IN_7 => UNWINDOWED_786 ,
										MUX_10_1_IN_8 => UNWINDOWED_531 ,
										MUX_10_1_IN_9 => UNWINDOWED_531 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_777
									);
MUX_REORD_UNIT_778 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_778 ,
										MUX_10_1_IN_1 => UNWINDOWED_777 ,
										MUX_10_1_IN_2 => UNWINDOWED_780 ,
										MUX_10_1_IN_3 => UNWINDOWED_773 ,
										MUX_10_1_IN_4 => UNWINDOWED_788 ,
										MUX_10_1_IN_5 => UNWINDOWED_788 ,
										MUX_10_1_IN_6 => UNWINDOWED_788 ,
										MUX_10_1_IN_7 => UNWINDOWED_788 ,
										MUX_10_1_IN_8 => UNWINDOWED_533 ,
										MUX_10_1_IN_9 => UNWINDOWED_533 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_778
									);
MUX_REORD_UNIT_779 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_779 ,
										MUX_10_1_IN_1 => UNWINDOWED_779 ,
										MUX_10_1_IN_2 => UNWINDOWED_782 ,
										MUX_10_1_IN_3 => UNWINDOWED_775 ,
										MUX_10_1_IN_4 => UNWINDOWED_790 ,
										MUX_10_1_IN_5 => UNWINDOWED_790 ,
										MUX_10_1_IN_6 => UNWINDOWED_790 ,
										MUX_10_1_IN_7 => UNWINDOWED_790 ,
										MUX_10_1_IN_8 => UNWINDOWED_535 ,
										MUX_10_1_IN_9 => UNWINDOWED_535 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_779
									);
MUX_REORD_UNIT_780 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_780 ,
										MUX_10_1_IN_1 => UNWINDOWED_780 ,
										MUX_10_1_IN_2 => UNWINDOWED_777 ,
										MUX_10_1_IN_3 => UNWINDOWED_777 ,
										MUX_10_1_IN_4 => UNWINDOWED_792 ,
										MUX_10_1_IN_5 => UNWINDOWED_792 ,
										MUX_10_1_IN_6 => UNWINDOWED_792 ,
										MUX_10_1_IN_7 => UNWINDOWED_792 ,
										MUX_10_1_IN_8 => UNWINDOWED_537 ,
										MUX_10_1_IN_9 => UNWINDOWED_537 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_780
									);
MUX_REORD_UNIT_781 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_781 ,
										MUX_10_1_IN_1 => UNWINDOWED_782 ,
										MUX_10_1_IN_2 => UNWINDOWED_779 ,
										MUX_10_1_IN_3 => UNWINDOWED_779 ,
										MUX_10_1_IN_4 => UNWINDOWED_794 ,
										MUX_10_1_IN_5 => UNWINDOWED_794 ,
										MUX_10_1_IN_6 => UNWINDOWED_794 ,
										MUX_10_1_IN_7 => UNWINDOWED_794 ,
										MUX_10_1_IN_8 => UNWINDOWED_539 ,
										MUX_10_1_IN_9 => UNWINDOWED_539 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_781
									);
MUX_REORD_UNIT_782 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_782 ,
										MUX_10_1_IN_1 => UNWINDOWED_781 ,
										MUX_10_1_IN_2 => UNWINDOWED_781 ,
										MUX_10_1_IN_3 => UNWINDOWED_781 ,
										MUX_10_1_IN_4 => UNWINDOWED_796 ,
										MUX_10_1_IN_5 => UNWINDOWED_796 ,
										MUX_10_1_IN_6 => UNWINDOWED_796 ,
										MUX_10_1_IN_7 => UNWINDOWED_796 ,
										MUX_10_1_IN_8 => UNWINDOWED_541 ,
										MUX_10_1_IN_9 => UNWINDOWED_541 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_782
									);
MUX_REORD_UNIT_783 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_783 ,
										MUX_10_1_IN_1 => UNWINDOWED_783 ,
										MUX_10_1_IN_2 => UNWINDOWED_783 ,
										MUX_10_1_IN_3 => UNWINDOWED_783 ,
										MUX_10_1_IN_4 => UNWINDOWED_798 ,
										MUX_10_1_IN_5 => UNWINDOWED_798 ,
										MUX_10_1_IN_6 => UNWINDOWED_798 ,
										MUX_10_1_IN_7 => UNWINDOWED_798 ,
										MUX_10_1_IN_8 => UNWINDOWED_543 ,
										MUX_10_1_IN_9 => UNWINDOWED_543 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_783
									);
MUX_REORD_UNIT_784 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_784 ,
										MUX_10_1_IN_1 => UNWINDOWED_784 ,
										MUX_10_1_IN_2 => UNWINDOWED_784 ,
										MUX_10_1_IN_3 => UNWINDOWED_784 ,
										MUX_10_1_IN_4 => UNWINDOWED_769 ,
										MUX_10_1_IN_5 => UNWINDOWED_800 ,
										MUX_10_1_IN_6 => UNWINDOWED_800 ,
										MUX_10_1_IN_7 => UNWINDOWED_800 ,
										MUX_10_1_IN_8 => UNWINDOWED_545 ,
										MUX_10_1_IN_9 => UNWINDOWED_545 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_784
									);
MUX_REORD_UNIT_785 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_785 ,
										MUX_10_1_IN_1 => UNWINDOWED_786 ,
										MUX_10_1_IN_2 => UNWINDOWED_786 ,
										MUX_10_1_IN_3 => UNWINDOWED_786 ,
										MUX_10_1_IN_4 => UNWINDOWED_771 ,
										MUX_10_1_IN_5 => UNWINDOWED_802 ,
										MUX_10_1_IN_6 => UNWINDOWED_802 ,
										MUX_10_1_IN_7 => UNWINDOWED_802 ,
										MUX_10_1_IN_8 => UNWINDOWED_547 ,
										MUX_10_1_IN_9 => UNWINDOWED_547 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_785
									);
MUX_REORD_UNIT_786 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_786 ,
										MUX_10_1_IN_1 => UNWINDOWED_785 ,
										MUX_10_1_IN_2 => UNWINDOWED_788 ,
										MUX_10_1_IN_3 => UNWINDOWED_788 ,
										MUX_10_1_IN_4 => UNWINDOWED_773 ,
										MUX_10_1_IN_5 => UNWINDOWED_804 ,
										MUX_10_1_IN_6 => UNWINDOWED_804 ,
										MUX_10_1_IN_7 => UNWINDOWED_804 ,
										MUX_10_1_IN_8 => UNWINDOWED_549 ,
										MUX_10_1_IN_9 => UNWINDOWED_549 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_786
									);
MUX_REORD_UNIT_787 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_787 ,
										MUX_10_1_IN_1 => UNWINDOWED_787 ,
										MUX_10_1_IN_2 => UNWINDOWED_790 ,
										MUX_10_1_IN_3 => UNWINDOWED_790 ,
										MUX_10_1_IN_4 => UNWINDOWED_775 ,
										MUX_10_1_IN_5 => UNWINDOWED_806 ,
										MUX_10_1_IN_6 => UNWINDOWED_806 ,
										MUX_10_1_IN_7 => UNWINDOWED_806 ,
										MUX_10_1_IN_8 => UNWINDOWED_551 ,
										MUX_10_1_IN_9 => UNWINDOWED_551 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_787
									);
MUX_REORD_UNIT_788 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_788 ,
										MUX_10_1_IN_1 => UNWINDOWED_788 ,
										MUX_10_1_IN_2 => UNWINDOWED_785 ,
										MUX_10_1_IN_3 => UNWINDOWED_792 ,
										MUX_10_1_IN_4 => UNWINDOWED_777 ,
										MUX_10_1_IN_5 => UNWINDOWED_808 ,
										MUX_10_1_IN_6 => UNWINDOWED_808 ,
										MUX_10_1_IN_7 => UNWINDOWED_808 ,
										MUX_10_1_IN_8 => UNWINDOWED_553 ,
										MUX_10_1_IN_9 => UNWINDOWED_553 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_788
									);
MUX_REORD_UNIT_789 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_789 ,
										MUX_10_1_IN_1 => UNWINDOWED_790 ,
										MUX_10_1_IN_2 => UNWINDOWED_787 ,
										MUX_10_1_IN_3 => UNWINDOWED_794 ,
										MUX_10_1_IN_4 => UNWINDOWED_779 ,
										MUX_10_1_IN_5 => UNWINDOWED_810 ,
										MUX_10_1_IN_6 => UNWINDOWED_810 ,
										MUX_10_1_IN_7 => UNWINDOWED_810 ,
										MUX_10_1_IN_8 => UNWINDOWED_555 ,
										MUX_10_1_IN_9 => UNWINDOWED_555 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_789
									);
MUX_REORD_UNIT_790 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_790 ,
										MUX_10_1_IN_1 => UNWINDOWED_789 ,
										MUX_10_1_IN_2 => UNWINDOWED_789 ,
										MUX_10_1_IN_3 => UNWINDOWED_796 ,
										MUX_10_1_IN_4 => UNWINDOWED_781 ,
										MUX_10_1_IN_5 => UNWINDOWED_812 ,
										MUX_10_1_IN_6 => UNWINDOWED_812 ,
										MUX_10_1_IN_7 => UNWINDOWED_812 ,
										MUX_10_1_IN_8 => UNWINDOWED_557 ,
										MUX_10_1_IN_9 => UNWINDOWED_557 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_790
									);
MUX_REORD_UNIT_791 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_791 ,
										MUX_10_1_IN_1 => UNWINDOWED_791 ,
										MUX_10_1_IN_2 => UNWINDOWED_791 ,
										MUX_10_1_IN_3 => UNWINDOWED_798 ,
										MUX_10_1_IN_4 => UNWINDOWED_783 ,
										MUX_10_1_IN_5 => UNWINDOWED_814 ,
										MUX_10_1_IN_6 => UNWINDOWED_814 ,
										MUX_10_1_IN_7 => UNWINDOWED_814 ,
										MUX_10_1_IN_8 => UNWINDOWED_559 ,
										MUX_10_1_IN_9 => UNWINDOWED_559 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_791
									);
MUX_REORD_UNIT_792 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_792 ,
										MUX_10_1_IN_1 => UNWINDOWED_792 ,
										MUX_10_1_IN_2 => UNWINDOWED_792 ,
										MUX_10_1_IN_3 => UNWINDOWED_785 ,
										MUX_10_1_IN_4 => UNWINDOWED_785 ,
										MUX_10_1_IN_5 => UNWINDOWED_816 ,
										MUX_10_1_IN_6 => UNWINDOWED_816 ,
										MUX_10_1_IN_7 => UNWINDOWED_816 ,
										MUX_10_1_IN_8 => UNWINDOWED_561 ,
										MUX_10_1_IN_9 => UNWINDOWED_561 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_792
									);
MUX_REORD_UNIT_793 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_793 ,
										MUX_10_1_IN_1 => UNWINDOWED_794 ,
										MUX_10_1_IN_2 => UNWINDOWED_794 ,
										MUX_10_1_IN_3 => UNWINDOWED_787 ,
										MUX_10_1_IN_4 => UNWINDOWED_787 ,
										MUX_10_1_IN_5 => UNWINDOWED_818 ,
										MUX_10_1_IN_6 => UNWINDOWED_818 ,
										MUX_10_1_IN_7 => UNWINDOWED_818 ,
										MUX_10_1_IN_8 => UNWINDOWED_563 ,
										MUX_10_1_IN_9 => UNWINDOWED_563 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_793
									);
MUX_REORD_UNIT_794 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_794 ,
										MUX_10_1_IN_1 => UNWINDOWED_793 ,
										MUX_10_1_IN_2 => UNWINDOWED_796 ,
										MUX_10_1_IN_3 => UNWINDOWED_789 ,
										MUX_10_1_IN_4 => UNWINDOWED_789 ,
										MUX_10_1_IN_5 => UNWINDOWED_820 ,
										MUX_10_1_IN_6 => UNWINDOWED_820 ,
										MUX_10_1_IN_7 => UNWINDOWED_820 ,
										MUX_10_1_IN_8 => UNWINDOWED_565 ,
										MUX_10_1_IN_9 => UNWINDOWED_565 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_794
									);
MUX_REORD_UNIT_795 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_795 ,
										MUX_10_1_IN_1 => UNWINDOWED_795 ,
										MUX_10_1_IN_2 => UNWINDOWED_798 ,
										MUX_10_1_IN_3 => UNWINDOWED_791 ,
										MUX_10_1_IN_4 => UNWINDOWED_791 ,
										MUX_10_1_IN_5 => UNWINDOWED_822 ,
										MUX_10_1_IN_6 => UNWINDOWED_822 ,
										MUX_10_1_IN_7 => UNWINDOWED_822 ,
										MUX_10_1_IN_8 => UNWINDOWED_567 ,
										MUX_10_1_IN_9 => UNWINDOWED_567 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_795
									);
MUX_REORD_UNIT_796 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_796 ,
										MUX_10_1_IN_1 => UNWINDOWED_796 ,
										MUX_10_1_IN_2 => UNWINDOWED_793 ,
										MUX_10_1_IN_3 => UNWINDOWED_793 ,
										MUX_10_1_IN_4 => UNWINDOWED_793 ,
										MUX_10_1_IN_5 => UNWINDOWED_824 ,
										MUX_10_1_IN_6 => UNWINDOWED_824 ,
										MUX_10_1_IN_7 => UNWINDOWED_824 ,
										MUX_10_1_IN_8 => UNWINDOWED_569 ,
										MUX_10_1_IN_9 => UNWINDOWED_569 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_796
									);
MUX_REORD_UNIT_797 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_797 ,
										MUX_10_1_IN_1 => UNWINDOWED_798 ,
										MUX_10_1_IN_2 => UNWINDOWED_795 ,
										MUX_10_1_IN_3 => UNWINDOWED_795 ,
										MUX_10_1_IN_4 => UNWINDOWED_795 ,
										MUX_10_1_IN_5 => UNWINDOWED_826 ,
										MUX_10_1_IN_6 => UNWINDOWED_826 ,
										MUX_10_1_IN_7 => UNWINDOWED_826 ,
										MUX_10_1_IN_8 => UNWINDOWED_571 ,
										MUX_10_1_IN_9 => UNWINDOWED_571 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_797
									);
MUX_REORD_UNIT_798 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_798 ,
										MUX_10_1_IN_1 => UNWINDOWED_797 ,
										MUX_10_1_IN_2 => UNWINDOWED_797 ,
										MUX_10_1_IN_3 => UNWINDOWED_797 ,
										MUX_10_1_IN_4 => UNWINDOWED_797 ,
										MUX_10_1_IN_5 => UNWINDOWED_828 ,
										MUX_10_1_IN_6 => UNWINDOWED_828 ,
										MUX_10_1_IN_7 => UNWINDOWED_828 ,
										MUX_10_1_IN_8 => UNWINDOWED_573 ,
										MUX_10_1_IN_9 => UNWINDOWED_573 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_798
									);
MUX_REORD_UNIT_799 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_799 ,
										MUX_10_1_IN_1 => UNWINDOWED_799 ,
										MUX_10_1_IN_2 => UNWINDOWED_799 ,
										MUX_10_1_IN_3 => UNWINDOWED_799 ,
										MUX_10_1_IN_4 => UNWINDOWED_799 ,
										MUX_10_1_IN_5 => UNWINDOWED_830 ,
										MUX_10_1_IN_6 => UNWINDOWED_830 ,
										MUX_10_1_IN_7 => UNWINDOWED_830 ,
										MUX_10_1_IN_8 => UNWINDOWED_575 ,
										MUX_10_1_IN_9 => UNWINDOWED_575 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_799
									);
MUX_REORD_UNIT_800 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_800 ,
										MUX_10_1_IN_1 => UNWINDOWED_800 ,
										MUX_10_1_IN_2 => UNWINDOWED_800 ,
										MUX_10_1_IN_3 => UNWINDOWED_800 ,
										MUX_10_1_IN_4 => UNWINDOWED_800 ,
										MUX_10_1_IN_5 => UNWINDOWED_769 ,
										MUX_10_1_IN_6 => UNWINDOWED_832 ,
										MUX_10_1_IN_7 => UNWINDOWED_832 ,
										MUX_10_1_IN_8 => UNWINDOWED_577 ,
										MUX_10_1_IN_9 => UNWINDOWED_577 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_800
									);
MUX_REORD_UNIT_801 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_801 ,
										MUX_10_1_IN_1 => UNWINDOWED_802 ,
										MUX_10_1_IN_2 => UNWINDOWED_802 ,
										MUX_10_1_IN_3 => UNWINDOWED_802 ,
										MUX_10_1_IN_4 => UNWINDOWED_802 ,
										MUX_10_1_IN_5 => UNWINDOWED_771 ,
										MUX_10_1_IN_6 => UNWINDOWED_834 ,
										MUX_10_1_IN_7 => UNWINDOWED_834 ,
										MUX_10_1_IN_8 => UNWINDOWED_579 ,
										MUX_10_1_IN_9 => UNWINDOWED_579 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_801
									);
MUX_REORD_UNIT_802 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_802 ,
										MUX_10_1_IN_1 => UNWINDOWED_801 ,
										MUX_10_1_IN_2 => UNWINDOWED_804 ,
										MUX_10_1_IN_3 => UNWINDOWED_804 ,
										MUX_10_1_IN_4 => UNWINDOWED_804 ,
										MUX_10_1_IN_5 => UNWINDOWED_773 ,
										MUX_10_1_IN_6 => UNWINDOWED_836 ,
										MUX_10_1_IN_7 => UNWINDOWED_836 ,
										MUX_10_1_IN_8 => UNWINDOWED_581 ,
										MUX_10_1_IN_9 => UNWINDOWED_581 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_802
									);
MUX_REORD_UNIT_803 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_803 ,
										MUX_10_1_IN_1 => UNWINDOWED_803 ,
										MUX_10_1_IN_2 => UNWINDOWED_806 ,
										MUX_10_1_IN_3 => UNWINDOWED_806 ,
										MUX_10_1_IN_4 => UNWINDOWED_806 ,
										MUX_10_1_IN_5 => UNWINDOWED_775 ,
										MUX_10_1_IN_6 => UNWINDOWED_838 ,
										MUX_10_1_IN_7 => UNWINDOWED_838 ,
										MUX_10_1_IN_8 => UNWINDOWED_583 ,
										MUX_10_1_IN_9 => UNWINDOWED_583 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_803
									);
MUX_REORD_UNIT_804 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_804 ,
										MUX_10_1_IN_1 => UNWINDOWED_804 ,
										MUX_10_1_IN_2 => UNWINDOWED_801 ,
										MUX_10_1_IN_3 => UNWINDOWED_808 ,
										MUX_10_1_IN_4 => UNWINDOWED_808 ,
										MUX_10_1_IN_5 => UNWINDOWED_777 ,
										MUX_10_1_IN_6 => UNWINDOWED_840 ,
										MUX_10_1_IN_7 => UNWINDOWED_840 ,
										MUX_10_1_IN_8 => UNWINDOWED_585 ,
										MUX_10_1_IN_9 => UNWINDOWED_585 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_804
									);
MUX_REORD_UNIT_805 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_805 ,
										MUX_10_1_IN_1 => UNWINDOWED_806 ,
										MUX_10_1_IN_2 => UNWINDOWED_803 ,
										MUX_10_1_IN_3 => UNWINDOWED_810 ,
										MUX_10_1_IN_4 => UNWINDOWED_810 ,
										MUX_10_1_IN_5 => UNWINDOWED_779 ,
										MUX_10_1_IN_6 => UNWINDOWED_842 ,
										MUX_10_1_IN_7 => UNWINDOWED_842 ,
										MUX_10_1_IN_8 => UNWINDOWED_587 ,
										MUX_10_1_IN_9 => UNWINDOWED_587 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_805
									);
MUX_REORD_UNIT_806 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_806 ,
										MUX_10_1_IN_1 => UNWINDOWED_805 ,
										MUX_10_1_IN_2 => UNWINDOWED_805 ,
										MUX_10_1_IN_3 => UNWINDOWED_812 ,
										MUX_10_1_IN_4 => UNWINDOWED_812 ,
										MUX_10_1_IN_5 => UNWINDOWED_781 ,
										MUX_10_1_IN_6 => UNWINDOWED_844 ,
										MUX_10_1_IN_7 => UNWINDOWED_844 ,
										MUX_10_1_IN_8 => UNWINDOWED_589 ,
										MUX_10_1_IN_9 => UNWINDOWED_589 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_806
									);
MUX_REORD_UNIT_807 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_807 ,
										MUX_10_1_IN_1 => UNWINDOWED_807 ,
										MUX_10_1_IN_2 => UNWINDOWED_807 ,
										MUX_10_1_IN_3 => UNWINDOWED_814 ,
										MUX_10_1_IN_4 => UNWINDOWED_814 ,
										MUX_10_1_IN_5 => UNWINDOWED_783 ,
										MUX_10_1_IN_6 => UNWINDOWED_846 ,
										MUX_10_1_IN_7 => UNWINDOWED_846 ,
										MUX_10_1_IN_8 => UNWINDOWED_591 ,
										MUX_10_1_IN_9 => UNWINDOWED_591 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_807
									);
MUX_REORD_UNIT_808 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_808 ,
										MUX_10_1_IN_1 => UNWINDOWED_808 ,
										MUX_10_1_IN_2 => UNWINDOWED_808 ,
										MUX_10_1_IN_3 => UNWINDOWED_801 ,
										MUX_10_1_IN_4 => UNWINDOWED_816 ,
										MUX_10_1_IN_5 => UNWINDOWED_785 ,
										MUX_10_1_IN_6 => UNWINDOWED_848 ,
										MUX_10_1_IN_7 => UNWINDOWED_848 ,
										MUX_10_1_IN_8 => UNWINDOWED_593 ,
										MUX_10_1_IN_9 => UNWINDOWED_593 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_808
									);
MUX_REORD_UNIT_809 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_809 ,
										MUX_10_1_IN_1 => UNWINDOWED_810 ,
										MUX_10_1_IN_2 => UNWINDOWED_810 ,
										MUX_10_1_IN_3 => UNWINDOWED_803 ,
										MUX_10_1_IN_4 => UNWINDOWED_818 ,
										MUX_10_1_IN_5 => UNWINDOWED_787 ,
										MUX_10_1_IN_6 => UNWINDOWED_850 ,
										MUX_10_1_IN_7 => UNWINDOWED_850 ,
										MUX_10_1_IN_8 => UNWINDOWED_595 ,
										MUX_10_1_IN_9 => UNWINDOWED_595 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_809
									);
MUX_REORD_UNIT_810 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_810 ,
										MUX_10_1_IN_1 => UNWINDOWED_809 ,
										MUX_10_1_IN_2 => UNWINDOWED_812 ,
										MUX_10_1_IN_3 => UNWINDOWED_805 ,
										MUX_10_1_IN_4 => UNWINDOWED_820 ,
										MUX_10_1_IN_5 => UNWINDOWED_789 ,
										MUX_10_1_IN_6 => UNWINDOWED_852 ,
										MUX_10_1_IN_7 => UNWINDOWED_852 ,
										MUX_10_1_IN_8 => UNWINDOWED_597 ,
										MUX_10_1_IN_9 => UNWINDOWED_597 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_810
									);
MUX_REORD_UNIT_811 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_811 ,
										MUX_10_1_IN_1 => UNWINDOWED_811 ,
										MUX_10_1_IN_2 => UNWINDOWED_814 ,
										MUX_10_1_IN_3 => UNWINDOWED_807 ,
										MUX_10_1_IN_4 => UNWINDOWED_822 ,
										MUX_10_1_IN_5 => UNWINDOWED_791 ,
										MUX_10_1_IN_6 => UNWINDOWED_854 ,
										MUX_10_1_IN_7 => UNWINDOWED_854 ,
										MUX_10_1_IN_8 => UNWINDOWED_599 ,
										MUX_10_1_IN_9 => UNWINDOWED_599 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_811
									);
MUX_REORD_UNIT_812 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_812 ,
										MUX_10_1_IN_1 => UNWINDOWED_812 ,
										MUX_10_1_IN_2 => UNWINDOWED_809 ,
										MUX_10_1_IN_3 => UNWINDOWED_809 ,
										MUX_10_1_IN_4 => UNWINDOWED_824 ,
										MUX_10_1_IN_5 => UNWINDOWED_793 ,
										MUX_10_1_IN_6 => UNWINDOWED_856 ,
										MUX_10_1_IN_7 => UNWINDOWED_856 ,
										MUX_10_1_IN_8 => UNWINDOWED_601 ,
										MUX_10_1_IN_9 => UNWINDOWED_601 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_812
									);
MUX_REORD_UNIT_813 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_813 ,
										MUX_10_1_IN_1 => UNWINDOWED_814 ,
										MUX_10_1_IN_2 => UNWINDOWED_811 ,
										MUX_10_1_IN_3 => UNWINDOWED_811 ,
										MUX_10_1_IN_4 => UNWINDOWED_826 ,
										MUX_10_1_IN_5 => UNWINDOWED_795 ,
										MUX_10_1_IN_6 => UNWINDOWED_858 ,
										MUX_10_1_IN_7 => UNWINDOWED_858 ,
										MUX_10_1_IN_8 => UNWINDOWED_603 ,
										MUX_10_1_IN_9 => UNWINDOWED_603 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_813
									);
MUX_REORD_UNIT_814 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_814 ,
										MUX_10_1_IN_1 => UNWINDOWED_813 ,
										MUX_10_1_IN_2 => UNWINDOWED_813 ,
										MUX_10_1_IN_3 => UNWINDOWED_813 ,
										MUX_10_1_IN_4 => UNWINDOWED_828 ,
										MUX_10_1_IN_5 => UNWINDOWED_797 ,
										MUX_10_1_IN_6 => UNWINDOWED_860 ,
										MUX_10_1_IN_7 => UNWINDOWED_860 ,
										MUX_10_1_IN_8 => UNWINDOWED_605 ,
										MUX_10_1_IN_9 => UNWINDOWED_605 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_814
									);
MUX_REORD_UNIT_815 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_815 ,
										MUX_10_1_IN_1 => UNWINDOWED_815 ,
										MUX_10_1_IN_2 => UNWINDOWED_815 ,
										MUX_10_1_IN_3 => UNWINDOWED_815 ,
										MUX_10_1_IN_4 => UNWINDOWED_830 ,
										MUX_10_1_IN_5 => UNWINDOWED_799 ,
										MUX_10_1_IN_6 => UNWINDOWED_862 ,
										MUX_10_1_IN_7 => UNWINDOWED_862 ,
										MUX_10_1_IN_8 => UNWINDOWED_607 ,
										MUX_10_1_IN_9 => UNWINDOWED_607 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_815
									);
MUX_REORD_UNIT_816 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_816 ,
										MUX_10_1_IN_1 => UNWINDOWED_816 ,
										MUX_10_1_IN_2 => UNWINDOWED_816 ,
										MUX_10_1_IN_3 => UNWINDOWED_816 ,
										MUX_10_1_IN_4 => UNWINDOWED_801 ,
										MUX_10_1_IN_5 => UNWINDOWED_801 ,
										MUX_10_1_IN_6 => UNWINDOWED_864 ,
										MUX_10_1_IN_7 => UNWINDOWED_864 ,
										MUX_10_1_IN_8 => UNWINDOWED_609 ,
										MUX_10_1_IN_9 => UNWINDOWED_609 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_816
									);
MUX_REORD_UNIT_817 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_817 ,
										MUX_10_1_IN_1 => UNWINDOWED_818 ,
										MUX_10_1_IN_2 => UNWINDOWED_818 ,
										MUX_10_1_IN_3 => UNWINDOWED_818 ,
										MUX_10_1_IN_4 => UNWINDOWED_803 ,
										MUX_10_1_IN_5 => UNWINDOWED_803 ,
										MUX_10_1_IN_6 => UNWINDOWED_866 ,
										MUX_10_1_IN_7 => UNWINDOWED_866 ,
										MUX_10_1_IN_8 => UNWINDOWED_611 ,
										MUX_10_1_IN_9 => UNWINDOWED_611 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_817
									);
MUX_REORD_UNIT_818 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_818 ,
										MUX_10_1_IN_1 => UNWINDOWED_817 ,
										MUX_10_1_IN_2 => UNWINDOWED_820 ,
										MUX_10_1_IN_3 => UNWINDOWED_820 ,
										MUX_10_1_IN_4 => UNWINDOWED_805 ,
										MUX_10_1_IN_5 => UNWINDOWED_805 ,
										MUX_10_1_IN_6 => UNWINDOWED_868 ,
										MUX_10_1_IN_7 => UNWINDOWED_868 ,
										MUX_10_1_IN_8 => UNWINDOWED_613 ,
										MUX_10_1_IN_9 => UNWINDOWED_613 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_818
									);
MUX_REORD_UNIT_819 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_819 ,
										MUX_10_1_IN_1 => UNWINDOWED_819 ,
										MUX_10_1_IN_2 => UNWINDOWED_822 ,
										MUX_10_1_IN_3 => UNWINDOWED_822 ,
										MUX_10_1_IN_4 => UNWINDOWED_807 ,
										MUX_10_1_IN_5 => UNWINDOWED_807 ,
										MUX_10_1_IN_6 => UNWINDOWED_870 ,
										MUX_10_1_IN_7 => UNWINDOWED_870 ,
										MUX_10_1_IN_8 => UNWINDOWED_615 ,
										MUX_10_1_IN_9 => UNWINDOWED_615 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_819
									);
MUX_REORD_UNIT_820 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_820 ,
										MUX_10_1_IN_1 => UNWINDOWED_820 ,
										MUX_10_1_IN_2 => UNWINDOWED_817 ,
										MUX_10_1_IN_3 => UNWINDOWED_824 ,
										MUX_10_1_IN_4 => UNWINDOWED_809 ,
										MUX_10_1_IN_5 => UNWINDOWED_809 ,
										MUX_10_1_IN_6 => UNWINDOWED_872 ,
										MUX_10_1_IN_7 => UNWINDOWED_872 ,
										MUX_10_1_IN_8 => UNWINDOWED_617 ,
										MUX_10_1_IN_9 => UNWINDOWED_617 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_820
									);
MUX_REORD_UNIT_821 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_821 ,
										MUX_10_1_IN_1 => UNWINDOWED_822 ,
										MUX_10_1_IN_2 => UNWINDOWED_819 ,
										MUX_10_1_IN_3 => UNWINDOWED_826 ,
										MUX_10_1_IN_4 => UNWINDOWED_811 ,
										MUX_10_1_IN_5 => UNWINDOWED_811 ,
										MUX_10_1_IN_6 => UNWINDOWED_874 ,
										MUX_10_1_IN_7 => UNWINDOWED_874 ,
										MUX_10_1_IN_8 => UNWINDOWED_619 ,
										MUX_10_1_IN_9 => UNWINDOWED_619 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_821
									);
MUX_REORD_UNIT_822 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_822 ,
										MUX_10_1_IN_1 => UNWINDOWED_821 ,
										MUX_10_1_IN_2 => UNWINDOWED_821 ,
										MUX_10_1_IN_3 => UNWINDOWED_828 ,
										MUX_10_1_IN_4 => UNWINDOWED_813 ,
										MUX_10_1_IN_5 => UNWINDOWED_813 ,
										MUX_10_1_IN_6 => UNWINDOWED_876 ,
										MUX_10_1_IN_7 => UNWINDOWED_876 ,
										MUX_10_1_IN_8 => UNWINDOWED_621 ,
										MUX_10_1_IN_9 => UNWINDOWED_621 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_822
									);
MUX_REORD_UNIT_823 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_823 ,
										MUX_10_1_IN_1 => UNWINDOWED_823 ,
										MUX_10_1_IN_2 => UNWINDOWED_823 ,
										MUX_10_1_IN_3 => UNWINDOWED_830 ,
										MUX_10_1_IN_4 => UNWINDOWED_815 ,
										MUX_10_1_IN_5 => UNWINDOWED_815 ,
										MUX_10_1_IN_6 => UNWINDOWED_878 ,
										MUX_10_1_IN_7 => UNWINDOWED_878 ,
										MUX_10_1_IN_8 => UNWINDOWED_623 ,
										MUX_10_1_IN_9 => UNWINDOWED_623 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_823
									);
MUX_REORD_UNIT_824 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_824 ,
										MUX_10_1_IN_1 => UNWINDOWED_824 ,
										MUX_10_1_IN_2 => UNWINDOWED_824 ,
										MUX_10_1_IN_3 => UNWINDOWED_817 ,
										MUX_10_1_IN_4 => UNWINDOWED_817 ,
										MUX_10_1_IN_5 => UNWINDOWED_817 ,
										MUX_10_1_IN_6 => UNWINDOWED_880 ,
										MUX_10_1_IN_7 => UNWINDOWED_880 ,
										MUX_10_1_IN_8 => UNWINDOWED_625 ,
										MUX_10_1_IN_9 => UNWINDOWED_625 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_824
									);
MUX_REORD_UNIT_825 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_825 ,
										MUX_10_1_IN_1 => UNWINDOWED_826 ,
										MUX_10_1_IN_2 => UNWINDOWED_826 ,
										MUX_10_1_IN_3 => UNWINDOWED_819 ,
										MUX_10_1_IN_4 => UNWINDOWED_819 ,
										MUX_10_1_IN_5 => UNWINDOWED_819 ,
										MUX_10_1_IN_6 => UNWINDOWED_882 ,
										MUX_10_1_IN_7 => UNWINDOWED_882 ,
										MUX_10_1_IN_8 => UNWINDOWED_627 ,
										MUX_10_1_IN_9 => UNWINDOWED_627 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_825
									);
MUX_REORD_UNIT_826 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_826 ,
										MUX_10_1_IN_1 => UNWINDOWED_825 ,
										MUX_10_1_IN_2 => UNWINDOWED_828 ,
										MUX_10_1_IN_3 => UNWINDOWED_821 ,
										MUX_10_1_IN_4 => UNWINDOWED_821 ,
										MUX_10_1_IN_5 => UNWINDOWED_821 ,
										MUX_10_1_IN_6 => UNWINDOWED_884 ,
										MUX_10_1_IN_7 => UNWINDOWED_884 ,
										MUX_10_1_IN_8 => UNWINDOWED_629 ,
										MUX_10_1_IN_9 => UNWINDOWED_629 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_826
									);
MUX_REORD_UNIT_827 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_827 ,
										MUX_10_1_IN_1 => UNWINDOWED_827 ,
										MUX_10_1_IN_2 => UNWINDOWED_830 ,
										MUX_10_1_IN_3 => UNWINDOWED_823 ,
										MUX_10_1_IN_4 => UNWINDOWED_823 ,
										MUX_10_1_IN_5 => UNWINDOWED_823 ,
										MUX_10_1_IN_6 => UNWINDOWED_886 ,
										MUX_10_1_IN_7 => UNWINDOWED_886 ,
										MUX_10_1_IN_8 => UNWINDOWED_631 ,
										MUX_10_1_IN_9 => UNWINDOWED_631 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_827
									);
MUX_REORD_UNIT_828 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_828 ,
										MUX_10_1_IN_1 => UNWINDOWED_828 ,
										MUX_10_1_IN_2 => UNWINDOWED_825 ,
										MUX_10_1_IN_3 => UNWINDOWED_825 ,
										MUX_10_1_IN_4 => UNWINDOWED_825 ,
										MUX_10_1_IN_5 => UNWINDOWED_825 ,
										MUX_10_1_IN_6 => UNWINDOWED_888 ,
										MUX_10_1_IN_7 => UNWINDOWED_888 ,
										MUX_10_1_IN_8 => UNWINDOWED_633 ,
										MUX_10_1_IN_9 => UNWINDOWED_633 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_828
									);
MUX_REORD_UNIT_829 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_829 ,
										MUX_10_1_IN_1 => UNWINDOWED_830 ,
										MUX_10_1_IN_2 => UNWINDOWED_827 ,
										MUX_10_1_IN_3 => UNWINDOWED_827 ,
										MUX_10_1_IN_4 => UNWINDOWED_827 ,
										MUX_10_1_IN_5 => UNWINDOWED_827 ,
										MUX_10_1_IN_6 => UNWINDOWED_890 ,
										MUX_10_1_IN_7 => UNWINDOWED_890 ,
										MUX_10_1_IN_8 => UNWINDOWED_635 ,
										MUX_10_1_IN_9 => UNWINDOWED_635 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_829
									);
MUX_REORD_UNIT_830 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_830 ,
										MUX_10_1_IN_1 => UNWINDOWED_829 ,
										MUX_10_1_IN_2 => UNWINDOWED_829 ,
										MUX_10_1_IN_3 => UNWINDOWED_829 ,
										MUX_10_1_IN_4 => UNWINDOWED_829 ,
										MUX_10_1_IN_5 => UNWINDOWED_829 ,
										MUX_10_1_IN_6 => UNWINDOWED_892 ,
										MUX_10_1_IN_7 => UNWINDOWED_892 ,
										MUX_10_1_IN_8 => UNWINDOWED_637 ,
										MUX_10_1_IN_9 => UNWINDOWED_637 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_830
									);
MUX_REORD_UNIT_831 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_831 ,
										MUX_10_1_IN_1 => UNWINDOWED_831 ,
										MUX_10_1_IN_2 => UNWINDOWED_831 ,
										MUX_10_1_IN_3 => UNWINDOWED_831 ,
										MUX_10_1_IN_4 => UNWINDOWED_831 ,
										MUX_10_1_IN_5 => UNWINDOWED_831 ,
										MUX_10_1_IN_6 => UNWINDOWED_894 ,
										MUX_10_1_IN_7 => UNWINDOWED_894 ,
										MUX_10_1_IN_8 => UNWINDOWED_639 ,
										MUX_10_1_IN_9 => UNWINDOWED_639 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_831
									);
MUX_REORD_UNIT_832 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_832 ,
										MUX_10_1_IN_1 => UNWINDOWED_832 ,
										MUX_10_1_IN_2 => UNWINDOWED_832 ,
										MUX_10_1_IN_3 => UNWINDOWED_832 ,
										MUX_10_1_IN_4 => UNWINDOWED_832 ,
										MUX_10_1_IN_5 => UNWINDOWED_832 ,
										MUX_10_1_IN_6 => UNWINDOWED_769 ,
										MUX_10_1_IN_7 => UNWINDOWED_896 ,
										MUX_10_1_IN_8 => UNWINDOWED_641 ,
										MUX_10_1_IN_9 => UNWINDOWED_641 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_832
									);
MUX_REORD_UNIT_833 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_833 ,
										MUX_10_1_IN_1 => UNWINDOWED_834 ,
										MUX_10_1_IN_2 => UNWINDOWED_834 ,
										MUX_10_1_IN_3 => UNWINDOWED_834 ,
										MUX_10_1_IN_4 => UNWINDOWED_834 ,
										MUX_10_1_IN_5 => UNWINDOWED_834 ,
										MUX_10_1_IN_6 => UNWINDOWED_771 ,
										MUX_10_1_IN_7 => UNWINDOWED_898 ,
										MUX_10_1_IN_8 => UNWINDOWED_643 ,
										MUX_10_1_IN_9 => UNWINDOWED_643 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_833
									);
MUX_REORD_UNIT_834 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_834 ,
										MUX_10_1_IN_1 => UNWINDOWED_833 ,
										MUX_10_1_IN_2 => UNWINDOWED_836 ,
										MUX_10_1_IN_3 => UNWINDOWED_836 ,
										MUX_10_1_IN_4 => UNWINDOWED_836 ,
										MUX_10_1_IN_5 => UNWINDOWED_836 ,
										MUX_10_1_IN_6 => UNWINDOWED_773 ,
										MUX_10_1_IN_7 => UNWINDOWED_900 ,
										MUX_10_1_IN_8 => UNWINDOWED_645 ,
										MUX_10_1_IN_9 => UNWINDOWED_645 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_834
									);
MUX_REORD_UNIT_835 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_835 ,
										MUX_10_1_IN_1 => UNWINDOWED_835 ,
										MUX_10_1_IN_2 => UNWINDOWED_838 ,
										MUX_10_1_IN_3 => UNWINDOWED_838 ,
										MUX_10_1_IN_4 => UNWINDOWED_838 ,
										MUX_10_1_IN_5 => UNWINDOWED_838 ,
										MUX_10_1_IN_6 => UNWINDOWED_775 ,
										MUX_10_1_IN_7 => UNWINDOWED_902 ,
										MUX_10_1_IN_8 => UNWINDOWED_647 ,
										MUX_10_1_IN_9 => UNWINDOWED_647 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_835
									);
MUX_REORD_UNIT_836 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_836 ,
										MUX_10_1_IN_1 => UNWINDOWED_836 ,
										MUX_10_1_IN_2 => UNWINDOWED_833 ,
										MUX_10_1_IN_3 => UNWINDOWED_840 ,
										MUX_10_1_IN_4 => UNWINDOWED_840 ,
										MUX_10_1_IN_5 => UNWINDOWED_840 ,
										MUX_10_1_IN_6 => UNWINDOWED_777 ,
										MUX_10_1_IN_7 => UNWINDOWED_904 ,
										MUX_10_1_IN_8 => UNWINDOWED_649 ,
										MUX_10_1_IN_9 => UNWINDOWED_649 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_836
									);
MUX_REORD_UNIT_837 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_837 ,
										MUX_10_1_IN_1 => UNWINDOWED_838 ,
										MUX_10_1_IN_2 => UNWINDOWED_835 ,
										MUX_10_1_IN_3 => UNWINDOWED_842 ,
										MUX_10_1_IN_4 => UNWINDOWED_842 ,
										MUX_10_1_IN_5 => UNWINDOWED_842 ,
										MUX_10_1_IN_6 => UNWINDOWED_779 ,
										MUX_10_1_IN_7 => UNWINDOWED_906 ,
										MUX_10_1_IN_8 => UNWINDOWED_651 ,
										MUX_10_1_IN_9 => UNWINDOWED_651 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_837
									);
MUX_REORD_UNIT_838 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_838 ,
										MUX_10_1_IN_1 => UNWINDOWED_837 ,
										MUX_10_1_IN_2 => UNWINDOWED_837 ,
										MUX_10_1_IN_3 => UNWINDOWED_844 ,
										MUX_10_1_IN_4 => UNWINDOWED_844 ,
										MUX_10_1_IN_5 => UNWINDOWED_844 ,
										MUX_10_1_IN_6 => UNWINDOWED_781 ,
										MUX_10_1_IN_7 => UNWINDOWED_908 ,
										MUX_10_1_IN_8 => UNWINDOWED_653 ,
										MUX_10_1_IN_9 => UNWINDOWED_653 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_838
									);
MUX_REORD_UNIT_839 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_839 ,
										MUX_10_1_IN_1 => UNWINDOWED_839 ,
										MUX_10_1_IN_2 => UNWINDOWED_839 ,
										MUX_10_1_IN_3 => UNWINDOWED_846 ,
										MUX_10_1_IN_4 => UNWINDOWED_846 ,
										MUX_10_1_IN_5 => UNWINDOWED_846 ,
										MUX_10_1_IN_6 => UNWINDOWED_783 ,
										MUX_10_1_IN_7 => UNWINDOWED_910 ,
										MUX_10_1_IN_8 => UNWINDOWED_655 ,
										MUX_10_1_IN_9 => UNWINDOWED_655 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_839
									);
MUX_REORD_UNIT_840 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_840 ,
										MUX_10_1_IN_1 => UNWINDOWED_840 ,
										MUX_10_1_IN_2 => UNWINDOWED_840 ,
										MUX_10_1_IN_3 => UNWINDOWED_833 ,
										MUX_10_1_IN_4 => UNWINDOWED_848 ,
										MUX_10_1_IN_5 => UNWINDOWED_848 ,
										MUX_10_1_IN_6 => UNWINDOWED_785 ,
										MUX_10_1_IN_7 => UNWINDOWED_912 ,
										MUX_10_1_IN_8 => UNWINDOWED_657 ,
										MUX_10_1_IN_9 => UNWINDOWED_657 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_840
									);
MUX_REORD_UNIT_841 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_841 ,
										MUX_10_1_IN_1 => UNWINDOWED_842 ,
										MUX_10_1_IN_2 => UNWINDOWED_842 ,
										MUX_10_1_IN_3 => UNWINDOWED_835 ,
										MUX_10_1_IN_4 => UNWINDOWED_850 ,
										MUX_10_1_IN_5 => UNWINDOWED_850 ,
										MUX_10_1_IN_6 => UNWINDOWED_787 ,
										MUX_10_1_IN_7 => UNWINDOWED_914 ,
										MUX_10_1_IN_8 => UNWINDOWED_659 ,
										MUX_10_1_IN_9 => UNWINDOWED_659 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_841
									);
MUX_REORD_UNIT_842 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_842 ,
										MUX_10_1_IN_1 => UNWINDOWED_841 ,
										MUX_10_1_IN_2 => UNWINDOWED_844 ,
										MUX_10_1_IN_3 => UNWINDOWED_837 ,
										MUX_10_1_IN_4 => UNWINDOWED_852 ,
										MUX_10_1_IN_5 => UNWINDOWED_852 ,
										MUX_10_1_IN_6 => UNWINDOWED_789 ,
										MUX_10_1_IN_7 => UNWINDOWED_916 ,
										MUX_10_1_IN_8 => UNWINDOWED_661 ,
										MUX_10_1_IN_9 => UNWINDOWED_661 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_842
									);
MUX_REORD_UNIT_843 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_843 ,
										MUX_10_1_IN_1 => UNWINDOWED_843 ,
										MUX_10_1_IN_2 => UNWINDOWED_846 ,
										MUX_10_1_IN_3 => UNWINDOWED_839 ,
										MUX_10_1_IN_4 => UNWINDOWED_854 ,
										MUX_10_1_IN_5 => UNWINDOWED_854 ,
										MUX_10_1_IN_6 => UNWINDOWED_791 ,
										MUX_10_1_IN_7 => UNWINDOWED_918 ,
										MUX_10_1_IN_8 => UNWINDOWED_663 ,
										MUX_10_1_IN_9 => UNWINDOWED_663 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_843
									);
MUX_REORD_UNIT_844 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_844 ,
										MUX_10_1_IN_1 => UNWINDOWED_844 ,
										MUX_10_1_IN_2 => UNWINDOWED_841 ,
										MUX_10_1_IN_3 => UNWINDOWED_841 ,
										MUX_10_1_IN_4 => UNWINDOWED_856 ,
										MUX_10_1_IN_5 => UNWINDOWED_856 ,
										MUX_10_1_IN_6 => UNWINDOWED_793 ,
										MUX_10_1_IN_7 => UNWINDOWED_920 ,
										MUX_10_1_IN_8 => UNWINDOWED_665 ,
										MUX_10_1_IN_9 => UNWINDOWED_665 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_844
									);
MUX_REORD_UNIT_845 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_845 ,
										MUX_10_1_IN_1 => UNWINDOWED_846 ,
										MUX_10_1_IN_2 => UNWINDOWED_843 ,
										MUX_10_1_IN_3 => UNWINDOWED_843 ,
										MUX_10_1_IN_4 => UNWINDOWED_858 ,
										MUX_10_1_IN_5 => UNWINDOWED_858 ,
										MUX_10_1_IN_6 => UNWINDOWED_795 ,
										MUX_10_1_IN_7 => UNWINDOWED_922 ,
										MUX_10_1_IN_8 => UNWINDOWED_667 ,
										MUX_10_1_IN_9 => UNWINDOWED_667 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_845
									);
MUX_REORD_UNIT_846 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_846 ,
										MUX_10_1_IN_1 => UNWINDOWED_845 ,
										MUX_10_1_IN_2 => UNWINDOWED_845 ,
										MUX_10_1_IN_3 => UNWINDOWED_845 ,
										MUX_10_1_IN_4 => UNWINDOWED_860 ,
										MUX_10_1_IN_5 => UNWINDOWED_860 ,
										MUX_10_1_IN_6 => UNWINDOWED_797 ,
										MUX_10_1_IN_7 => UNWINDOWED_924 ,
										MUX_10_1_IN_8 => UNWINDOWED_669 ,
										MUX_10_1_IN_9 => UNWINDOWED_669 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_846
									);
MUX_REORD_UNIT_847 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_847 ,
										MUX_10_1_IN_1 => UNWINDOWED_847 ,
										MUX_10_1_IN_2 => UNWINDOWED_847 ,
										MUX_10_1_IN_3 => UNWINDOWED_847 ,
										MUX_10_1_IN_4 => UNWINDOWED_862 ,
										MUX_10_1_IN_5 => UNWINDOWED_862 ,
										MUX_10_1_IN_6 => UNWINDOWED_799 ,
										MUX_10_1_IN_7 => UNWINDOWED_926 ,
										MUX_10_1_IN_8 => UNWINDOWED_671 ,
										MUX_10_1_IN_9 => UNWINDOWED_671 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_847
									);
MUX_REORD_UNIT_848 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_848 ,
										MUX_10_1_IN_1 => UNWINDOWED_848 ,
										MUX_10_1_IN_2 => UNWINDOWED_848 ,
										MUX_10_1_IN_3 => UNWINDOWED_848 ,
										MUX_10_1_IN_4 => UNWINDOWED_833 ,
										MUX_10_1_IN_5 => UNWINDOWED_864 ,
										MUX_10_1_IN_6 => UNWINDOWED_801 ,
										MUX_10_1_IN_7 => UNWINDOWED_928 ,
										MUX_10_1_IN_8 => UNWINDOWED_673 ,
										MUX_10_1_IN_9 => UNWINDOWED_673 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_848
									);
MUX_REORD_UNIT_849 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_849 ,
										MUX_10_1_IN_1 => UNWINDOWED_850 ,
										MUX_10_1_IN_2 => UNWINDOWED_850 ,
										MUX_10_1_IN_3 => UNWINDOWED_850 ,
										MUX_10_1_IN_4 => UNWINDOWED_835 ,
										MUX_10_1_IN_5 => UNWINDOWED_866 ,
										MUX_10_1_IN_6 => UNWINDOWED_803 ,
										MUX_10_1_IN_7 => UNWINDOWED_930 ,
										MUX_10_1_IN_8 => UNWINDOWED_675 ,
										MUX_10_1_IN_9 => UNWINDOWED_675 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_849
									);
MUX_REORD_UNIT_850 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_850 ,
										MUX_10_1_IN_1 => UNWINDOWED_849 ,
										MUX_10_1_IN_2 => UNWINDOWED_852 ,
										MUX_10_1_IN_3 => UNWINDOWED_852 ,
										MUX_10_1_IN_4 => UNWINDOWED_837 ,
										MUX_10_1_IN_5 => UNWINDOWED_868 ,
										MUX_10_1_IN_6 => UNWINDOWED_805 ,
										MUX_10_1_IN_7 => UNWINDOWED_932 ,
										MUX_10_1_IN_8 => UNWINDOWED_677 ,
										MUX_10_1_IN_9 => UNWINDOWED_677 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_850
									);
MUX_REORD_UNIT_851 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_851 ,
										MUX_10_1_IN_1 => UNWINDOWED_851 ,
										MUX_10_1_IN_2 => UNWINDOWED_854 ,
										MUX_10_1_IN_3 => UNWINDOWED_854 ,
										MUX_10_1_IN_4 => UNWINDOWED_839 ,
										MUX_10_1_IN_5 => UNWINDOWED_870 ,
										MUX_10_1_IN_6 => UNWINDOWED_807 ,
										MUX_10_1_IN_7 => UNWINDOWED_934 ,
										MUX_10_1_IN_8 => UNWINDOWED_679 ,
										MUX_10_1_IN_9 => UNWINDOWED_679 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_851
									);
MUX_REORD_UNIT_852 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_852 ,
										MUX_10_1_IN_1 => UNWINDOWED_852 ,
										MUX_10_1_IN_2 => UNWINDOWED_849 ,
										MUX_10_1_IN_3 => UNWINDOWED_856 ,
										MUX_10_1_IN_4 => UNWINDOWED_841 ,
										MUX_10_1_IN_5 => UNWINDOWED_872 ,
										MUX_10_1_IN_6 => UNWINDOWED_809 ,
										MUX_10_1_IN_7 => UNWINDOWED_936 ,
										MUX_10_1_IN_8 => UNWINDOWED_681 ,
										MUX_10_1_IN_9 => UNWINDOWED_681 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_852
									);
MUX_REORD_UNIT_853 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_853 ,
										MUX_10_1_IN_1 => UNWINDOWED_854 ,
										MUX_10_1_IN_2 => UNWINDOWED_851 ,
										MUX_10_1_IN_3 => UNWINDOWED_858 ,
										MUX_10_1_IN_4 => UNWINDOWED_843 ,
										MUX_10_1_IN_5 => UNWINDOWED_874 ,
										MUX_10_1_IN_6 => UNWINDOWED_811 ,
										MUX_10_1_IN_7 => UNWINDOWED_938 ,
										MUX_10_1_IN_8 => UNWINDOWED_683 ,
										MUX_10_1_IN_9 => UNWINDOWED_683 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_853
									);
MUX_REORD_UNIT_854 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_854 ,
										MUX_10_1_IN_1 => UNWINDOWED_853 ,
										MUX_10_1_IN_2 => UNWINDOWED_853 ,
										MUX_10_1_IN_3 => UNWINDOWED_860 ,
										MUX_10_1_IN_4 => UNWINDOWED_845 ,
										MUX_10_1_IN_5 => UNWINDOWED_876 ,
										MUX_10_1_IN_6 => UNWINDOWED_813 ,
										MUX_10_1_IN_7 => UNWINDOWED_940 ,
										MUX_10_1_IN_8 => UNWINDOWED_685 ,
										MUX_10_1_IN_9 => UNWINDOWED_685 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_854
									);
MUX_REORD_UNIT_855 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_855 ,
										MUX_10_1_IN_1 => UNWINDOWED_855 ,
										MUX_10_1_IN_2 => UNWINDOWED_855 ,
										MUX_10_1_IN_3 => UNWINDOWED_862 ,
										MUX_10_1_IN_4 => UNWINDOWED_847 ,
										MUX_10_1_IN_5 => UNWINDOWED_878 ,
										MUX_10_1_IN_6 => UNWINDOWED_815 ,
										MUX_10_1_IN_7 => UNWINDOWED_942 ,
										MUX_10_1_IN_8 => UNWINDOWED_687 ,
										MUX_10_1_IN_9 => UNWINDOWED_687 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_855
									);
MUX_REORD_UNIT_856 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_856 ,
										MUX_10_1_IN_1 => UNWINDOWED_856 ,
										MUX_10_1_IN_2 => UNWINDOWED_856 ,
										MUX_10_1_IN_3 => UNWINDOWED_849 ,
										MUX_10_1_IN_4 => UNWINDOWED_849 ,
										MUX_10_1_IN_5 => UNWINDOWED_880 ,
										MUX_10_1_IN_6 => UNWINDOWED_817 ,
										MUX_10_1_IN_7 => UNWINDOWED_944 ,
										MUX_10_1_IN_8 => UNWINDOWED_689 ,
										MUX_10_1_IN_9 => UNWINDOWED_689 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_856
									);
MUX_REORD_UNIT_857 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_857 ,
										MUX_10_1_IN_1 => UNWINDOWED_858 ,
										MUX_10_1_IN_2 => UNWINDOWED_858 ,
										MUX_10_1_IN_3 => UNWINDOWED_851 ,
										MUX_10_1_IN_4 => UNWINDOWED_851 ,
										MUX_10_1_IN_5 => UNWINDOWED_882 ,
										MUX_10_1_IN_6 => UNWINDOWED_819 ,
										MUX_10_1_IN_7 => UNWINDOWED_946 ,
										MUX_10_1_IN_8 => UNWINDOWED_691 ,
										MUX_10_1_IN_9 => UNWINDOWED_691 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_857
									);
MUX_REORD_UNIT_858 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_858 ,
										MUX_10_1_IN_1 => UNWINDOWED_857 ,
										MUX_10_1_IN_2 => UNWINDOWED_860 ,
										MUX_10_1_IN_3 => UNWINDOWED_853 ,
										MUX_10_1_IN_4 => UNWINDOWED_853 ,
										MUX_10_1_IN_5 => UNWINDOWED_884 ,
										MUX_10_1_IN_6 => UNWINDOWED_821 ,
										MUX_10_1_IN_7 => UNWINDOWED_948 ,
										MUX_10_1_IN_8 => UNWINDOWED_693 ,
										MUX_10_1_IN_9 => UNWINDOWED_693 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_858
									);
MUX_REORD_UNIT_859 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_859 ,
										MUX_10_1_IN_1 => UNWINDOWED_859 ,
										MUX_10_1_IN_2 => UNWINDOWED_862 ,
										MUX_10_1_IN_3 => UNWINDOWED_855 ,
										MUX_10_1_IN_4 => UNWINDOWED_855 ,
										MUX_10_1_IN_5 => UNWINDOWED_886 ,
										MUX_10_1_IN_6 => UNWINDOWED_823 ,
										MUX_10_1_IN_7 => UNWINDOWED_950 ,
										MUX_10_1_IN_8 => UNWINDOWED_695 ,
										MUX_10_1_IN_9 => UNWINDOWED_695 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_859
									);
MUX_REORD_UNIT_860 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_860 ,
										MUX_10_1_IN_1 => UNWINDOWED_860 ,
										MUX_10_1_IN_2 => UNWINDOWED_857 ,
										MUX_10_1_IN_3 => UNWINDOWED_857 ,
										MUX_10_1_IN_4 => UNWINDOWED_857 ,
										MUX_10_1_IN_5 => UNWINDOWED_888 ,
										MUX_10_1_IN_6 => UNWINDOWED_825 ,
										MUX_10_1_IN_7 => UNWINDOWED_952 ,
										MUX_10_1_IN_8 => UNWINDOWED_697 ,
										MUX_10_1_IN_9 => UNWINDOWED_697 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_860
									);
MUX_REORD_UNIT_861 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_861 ,
										MUX_10_1_IN_1 => UNWINDOWED_862 ,
										MUX_10_1_IN_2 => UNWINDOWED_859 ,
										MUX_10_1_IN_3 => UNWINDOWED_859 ,
										MUX_10_1_IN_4 => UNWINDOWED_859 ,
										MUX_10_1_IN_5 => UNWINDOWED_890 ,
										MUX_10_1_IN_6 => UNWINDOWED_827 ,
										MUX_10_1_IN_7 => UNWINDOWED_954 ,
										MUX_10_1_IN_8 => UNWINDOWED_699 ,
										MUX_10_1_IN_9 => UNWINDOWED_699 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_861
									);
MUX_REORD_UNIT_862 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_862 ,
										MUX_10_1_IN_1 => UNWINDOWED_861 ,
										MUX_10_1_IN_2 => UNWINDOWED_861 ,
										MUX_10_1_IN_3 => UNWINDOWED_861 ,
										MUX_10_1_IN_4 => UNWINDOWED_861 ,
										MUX_10_1_IN_5 => UNWINDOWED_892 ,
										MUX_10_1_IN_6 => UNWINDOWED_829 ,
										MUX_10_1_IN_7 => UNWINDOWED_956 ,
										MUX_10_1_IN_8 => UNWINDOWED_701 ,
										MUX_10_1_IN_9 => UNWINDOWED_701 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_862
									);
MUX_REORD_UNIT_863 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_863 ,
										MUX_10_1_IN_1 => UNWINDOWED_863 ,
										MUX_10_1_IN_2 => UNWINDOWED_863 ,
										MUX_10_1_IN_3 => UNWINDOWED_863 ,
										MUX_10_1_IN_4 => UNWINDOWED_863 ,
										MUX_10_1_IN_5 => UNWINDOWED_894 ,
										MUX_10_1_IN_6 => UNWINDOWED_831 ,
										MUX_10_1_IN_7 => UNWINDOWED_958 ,
										MUX_10_1_IN_8 => UNWINDOWED_703 ,
										MUX_10_1_IN_9 => UNWINDOWED_703 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_863
									);
MUX_REORD_UNIT_864 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_864 ,
										MUX_10_1_IN_1 => UNWINDOWED_864 ,
										MUX_10_1_IN_2 => UNWINDOWED_864 ,
										MUX_10_1_IN_3 => UNWINDOWED_864 ,
										MUX_10_1_IN_4 => UNWINDOWED_864 ,
										MUX_10_1_IN_5 => UNWINDOWED_833 ,
										MUX_10_1_IN_6 => UNWINDOWED_833 ,
										MUX_10_1_IN_7 => UNWINDOWED_960 ,
										MUX_10_1_IN_8 => UNWINDOWED_705 ,
										MUX_10_1_IN_9 => UNWINDOWED_705 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_864
									);
MUX_REORD_UNIT_865 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_865 ,
										MUX_10_1_IN_1 => UNWINDOWED_866 ,
										MUX_10_1_IN_2 => UNWINDOWED_866 ,
										MUX_10_1_IN_3 => UNWINDOWED_866 ,
										MUX_10_1_IN_4 => UNWINDOWED_866 ,
										MUX_10_1_IN_5 => UNWINDOWED_835 ,
										MUX_10_1_IN_6 => UNWINDOWED_835 ,
										MUX_10_1_IN_7 => UNWINDOWED_962 ,
										MUX_10_1_IN_8 => UNWINDOWED_707 ,
										MUX_10_1_IN_9 => UNWINDOWED_707 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_865
									);
MUX_REORD_UNIT_866 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_866 ,
										MUX_10_1_IN_1 => UNWINDOWED_865 ,
										MUX_10_1_IN_2 => UNWINDOWED_868 ,
										MUX_10_1_IN_3 => UNWINDOWED_868 ,
										MUX_10_1_IN_4 => UNWINDOWED_868 ,
										MUX_10_1_IN_5 => UNWINDOWED_837 ,
										MUX_10_1_IN_6 => UNWINDOWED_837 ,
										MUX_10_1_IN_7 => UNWINDOWED_964 ,
										MUX_10_1_IN_8 => UNWINDOWED_709 ,
										MUX_10_1_IN_9 => UNWINDOWED_709 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_866
									);
MUX_REORD_UNIT_867 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_867 ,
										MUX_10_1_IN_1 => UNWINDOWED_867 ,
										MUX_10_1_IN_2 => UNWINDOWED_870 ,
										MUX_10_1_IN_3 => UNWINDOWED_870 ,
										MUX_10_1_IN_4 => UNWINDOWED_870 ,
										MUX_10_1_IN_5 => UNWINDOWED_839 ,
										MUX_10_1_IN_6 => UNWINDOWED_839 ,
										MUX_10_1_IN_7 => UNWINDOWED_966 ,
										MUX_10_1_IN_8 => UNWINDOWED_711 ,
										MUX_10_1_IN_9 => UNWINDOWED_711 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_867
									);
MUX_REORD_UNIT_868 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_868 ,
										MUX_10_1_IN_1 => UNWINDOWED_868 ,
										MUX_10_1_IN_2 => UNWINDOWED_865 ,
										MUX_10_1_IN_3 => UNWINDOWED_872 ,
										MUX_10_1_IN_4 => UNWINDOWED_872 ,
										MUX_10_1_IN_5 => UNWINDOWED_841 ,
										MUX_10_1_IN_6 => UNWINDOWED_841 ,
										MUX_10_1_IN_7 => UNWINDOWED_968 ,
										MUX_10_1_IN_8 => UNWINDOWED_713 ,
										MUX_10_1_IN_9 => UNWINDOWED_713 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_868
									);
MUX_REORD_UNIT_869 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_869 ,
										MUX_10_1_IN_1 => UNWINDOWED_870 ,
										MUX_10_1_IN_2 => UNWINDOWED_867 ,
										MUX_10_1_IN_3 => UNWINDOWED_874 ,
										MUX_10_1_IN_4 => UNWINDOWED_874 ,
										MUX_10_1_IN_5 => UNWINDOWED_843 ,
										MUX_10_1_IN_6 => UNWINDOWED_843 ,
										MUX_10_1_IN_7 => UNWINDOWED_970 ,
										MUX_10_1_IN_8 => UNWINDOWED_715 ,
										MUX_10_1_IN_9 => UNWINDOWED_715 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_869
									);
MUX_REORD_UNIT_870 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_870 ,
										MUX_10_1_IN_1 => UNWINDOWED_869 ,
										MUX_10_1_IN_2 => UNWINDOWED_869 ,
										MUX_10_1_IN_3 => UNWINDOWED_876 ,
										MUX_10_1_IN_4 => UNWINDOWED_876 ,
										MUX_10_1_IN_5 => UNWINDOWED_845 ,
										MUX_10_1_IN_6 => UNWINDOWED_845 ,
										MUX_10_1_IN_7 => UNWINDOWED_972 ,
										MUX_10_1_IN_8 => UNWINDOWED_717 ,
										MUX_10_1_IN_9 => UNWINDOWED_717 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_870
									);
MUX_REORD_UNIT_871 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_871 ,
										MUX_10_1_IN_1 => UNWINDOWED_871 ,
										MUX_10_1_IN_2 => UNWINDOWED_871 ,
										MUX_10_1_IN_3 => UNWINDOWED_878 ,
										MUX_10_1_IN_4 => UNWINDOWED_878 ,
										MUX_10_1_IN_5 => UNWINDOWED_847 ,
										MUX_10_1_IN_6 => UNWINDOWED_847 ,
										MUX_10_1_IN_7 => UNWINDOWED_974 ,
										MUX_10_1_IN_8 => UNWINDOWED_719 ,
										MUX_10_1_IN_9 => UNWINDOWED_719 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_871
									);
MUX_REORD_UNIT_872 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_872 ,
										MUX_10_1_IN_1 => UNWINDOWED_872 ,
										MUX_10_1_IN_2 => UNWINDOWED_872 ,
										MUX_10_1_IN_3 => UNWINDOWED_865 ,
										MUX_10_1_IN_4 => UNWINDOWED_880 ,
										MUX_10_1_IN_5 => UNWINDOWED_849 ,
										MUX_10_1_IN_6 => UNWINDOWED_849 ,
										MUX_10_1_IN_7 => UNWINDOWED_976 ,
										MUX_10_1_IN_8 => UNWINDOWED_721 ,
										MUX_10_1_IN_9 => UNWINDOWED_721 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_872
									);
MUX_REORD_UNIT_873 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_873 ,
										MUX_10_1_IN_1 => UNWINDOWED_874 ,
										MUX_10_1_IN_2 => UNWINDOWED_874 ,
										MUX_10_1_IN_3 => UNWINDOWED_867 ,
										MUX_10_1_IN_4 => UNWINDOWED_882 ,
										MUX_10_1_IN_5 => UNWINDOWED_851 ,
										MUX_10_1_IN_6 => UNWINDOWED_851 ,
										MUX_10_1_IN_7 => UNWINDOWED_978 ,
										MUX_10_1_IN_8 => UNWINDOWED_723 ,
										MUX_10_1_IN_9 => UNWINDOWED_723 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_873
									);
MUX_REORD_UNIT_874 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_874 ,
										MUX_10_1_IN_1 => UNWINDOWED_873 ,
										MUX_10_1_IN_2 => UNWINDOWED_876 ,
										MUX_10_1_IN_3 => UNWINDOWED_869 ,
										MUX_10_1_IN_4 => UNWINDOWED_884 ,
										MUX_10_1_IN_5 => UNWINDOWED_853 ,
										MUX_10_1_IN_6 => UNWINDOWED_853 ,
										MUX_10_1_IN_7 => UNWINDOWED_980 ,
										MUX_10_1_IN_8 => UNWINDOWED_725 ,
										MUX_10_1_IN_9 => UNWINDOWED_725 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_874
									);
MUX_REORD_UNIT_875 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_875 ,
										MUX_10_1_IN_1 => UNWINDOWED_875 ,
										MUX_10_1_IN_2 => UNWINDOWED_878 ,
										MUX_10_1_IN_3 => UNWINDOWED_871 ,
										MUX_10_1_IN_4 => UNWINDOWED_886 ,
										MUX_10_1_IN_5 => UNWINDOWED_855 ,
										MUX_10_1_IN_6 => UNWINDOWED_855 ,
										MUX_10_1_IN_7 => UNWINDOWED_982 ,
										MUX_10_1_IN_8 => UNWINDOWED_727 ,
										MUX_10_1_IN_9 => UNWINDOWED_727 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_875
									);
MUX_REORD_UNIT_876 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_876 ,
										MUX_10_1_IN_1 => UNWINDOWED_876 ,
										MUX_10_1_IN_2 => UNWINDOWED_873 ,
										MUX_10_1_IN_3 => UNWINDOWED_873 ,
										MUX_10_1_IN_4 => UNWINDOWED_888 ,
										MUX_10_1_IN_5 => UNWINDOWED_857 ,
										MUX_10_1_IN_6 => UNWINDOWED_857 ,
										MUX_10_1_IN_7 => UNWINDOWED_984 ,
										MUX_10_1_IN_8 => UNWINDOWED_729 ,
										MUX_10_1_IN_9 => UNWINDOWED_729 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_876
									);
MUX_REORD_UNIT_877 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_877 ,
										MUX_10_1_IN_1 => UNWINDOWED_878 ,
										MUX_10_1_IN_2 => UNWINDOWED_875 ,
										MUX_10_1_IN_3 => UNWINDOWED_875 ,
										MUX_10_1_IN_4 => UNWINDOWED_890 ,
										MUX_10_1_IN_5 => UNWINDOWED_859 ,
										MUX_10_1_IN_6 => UNWINDOWED_859 ,
										MUX_10_1_IN_7 => UNWINDOWED_986 ,
										MUX_10_1_IN_8 => UNWINDOWED_731 ,
										MUX_10_1_IN_9 => UNWINDOWED_731 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_877
									);
MUX_REORD_UNIT_878 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_878 ,
										MUX_10_1_IN_1 => UNWINDOWED_877 ,
										MUX_10_1_IN_2 => UNWINDOWED_877 ,
										MUX_10_1_IN_3 => UNWINDOWED_877 ,
										MUX_10_1_IN_4 => UNWINDOWED_892 ,
										MUX_10_1_IN_5 => UNWINDOWED_861 ,
										MUX_10_1_IN_6 => UNWINDOWED_861 ,
										MUX_10_1_IN_7 => UNWINDOWED_988 ,
										MUX_10_1_IN_8 => UNWINDOWED_733 ,
										MUX_10_1_IN_9 => UNWINDOWED_733 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_878
									);
MUX_REORD_UNIT_879 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_879 ,
										MUX_10_1_IN_1 => UNWINDOWED_879 ,
										MUX_10_1_IN_2 => UNWINDOWED_879 ,
										MUX_10_1_IN_3 => UNWINDOWED_879 ,
										MUX_10_1_IN_4 => UNWINDOWED_894 ,
										MUX_10_1_IN_5 => UNWINDOWED_863 ,
										MUX_10_1_IN_6 => UNWINDOWED_863 ,
										MUX_10_1_IN_7 => UNWINDOWED_990 ,
										MUX_10_1_IN_8 => UNWINDOWED_735 ,
										MUX_10_1_IN_9 => UNWINDOWED_735 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_879
									);
MUX_REORD_UNIT_880 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_880 ,
										MUX_10_1_IN_1 => UNWINDOWED_880 ,
										MUX_10_1_IN_2 => UNWINDOWED_880 ,
										MUX_10_1_IN_3 => UNWINDOWED_880 ,
										MUX_10_1_IN_4 => UNWINDOWED_865 ,
										MUX_10_1_IN_5 => UNWINDOWED_865 ,
										MUX_10_1_IN_6 => UNWINDOWED_865 ,
										MUX_10_1_IN_7 => UNWINDOWED_992 ,
										MUX_10_1_IN_8 => UNWINDOWED_737 ,
										MUX_10_1_IN_9 => UNWINDOWED_737 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_880
									);
MUX_REORD_UNIT_881 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_881 ,
										MUX_10_1_IN_1 => UNWINDOWED_882 ,
										MUX_10_1_IN_2 => UNWINDOWED_882 ,
										MUX_10_1_IN_3 => UNWINDOWED_882 ,
										MUX_10_1_IN_4 => UNWINDOWED_867 ,
										MUX_10_1_IN_5 => UNWINDOWED_867 ,
										MUX_10_1_IN_6 => UNWINDOWED_867 ,
										MUX_10_1_IN_7 => UNWINDOWED_994 ,
										MUX_10_1_IN_8 => UNWINDOWED_739 ,
										MUX_10_1_IN_9 => UNWINDOWED_739 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_881
									);
MUX_REORD_UNIT_882 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_882 ,
										MUX_10_1_IN_1 => UNWINDOWED_881 ,
										MUX_10_1_IN_2 => UNWINDOWED_884 ,
										MUX_10_1_IN_3 => UNWINDOWED_884 ,
										MUX_10_1_IN_4 => UNWINDOWED_869 ,
										MUX_10_1_IN_5 => UNWINDOWED_869 ,
										MUX_10_1_IN_6 => UNWINDOWED_869 ,
										MUX_10_1_IN_7 => UNWINDOWED_996 ,
										MUX_10_1_IN_8 => UNWINDOWED_741 ,
										MUX_10_1_IN_9 => UNWINDOWED_741 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_882
									);
MUX_REORD_UNIT_883 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_883 ,
										MUX_10_1_IN_1 => UNWINDOWED_883 ,
										MUX_10_1_IN_2 => UNWINDOWED_886 ,
										MUX_10_1_IN_3 => UNWINDOWED_886 ,
										MUX_10_1_IN_4 => UNWINDOWED_871 ,
										MUX_10_1_IN_5 => UNWINDOWED_871 ,
										MUX_10_1_IN_6 => UNWINDOWED_871 ,
										MUX_10_1_IN_7 => UNWINDOWED_998 ,
										MUX_10_1_IN_8 => UNWINDOWED_743 ,
										MUX_10_1_IN_9 => UNWINDOWED_743 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_883
									);
MUX_REORD_UNIT_884 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_884 ,
										MUX_10_1_IN_1 => UNWINDOWED_884 ,
										MUX_10_1_IN_2 => UNWINDOWED_881 ,
										MUX_10_1_IN_3 => UNWINDOWED_888 ,
										MUX_10_1_IN_4 => UNWINDOWED_873 ,
										MUX_10_1_IN_5 => UNWINDOWED_873 ,
										MUX_10_1_IN_6 => UNWINDOWED_873 ,
										MUX_10_1_IN_7 => UNWINDOWED_1000 ,
										MUX_10_1_IN_8 => UNWINDOWED_745 ,
										MUX_10_1_IN_9 => UNWINDOWED_745 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_884
									);
MUX_REORD_UNIT_885 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_885 ,
										MUX_10_1_IN_1 => UNWINDOWED_886 ,
										MUX_10_1_IN_2 => UNWINDOWED_883 ,
										MUX_10_1_IN_3 => UNWINDOWED_890 ,
										MUX_10_1_IN_4 => UNWINDOWED_875 ,
										MUX_10_1_IN_5 => UNWINDOWED_875 ,
										MUX_10_1_IN_6 => UNWINDOWED_875 ,
										MUX_10_1_IN_7 => UNWINDOWED_1002 ,
										MUX_10_1_IN_8 => UNWINDOWED_747 ,
										MUX_10_1_IN_9 => UNWINDOWED_747 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_885
									);
MUX_REORD_UNIT_886 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_886 ,
										MUX_10_1_IN_1 => UNWINDOWED_885 ,
										MUX_10_1_IN_2 => UNWINDOWED_885 ,
										MUX_10_1_IN_3 => UNWINDOWED_892 ,
										MUX_10_1_IN_4 => UNWINDOWED_877 ,
										MUX_10_1_IN_5 => UNWINDOWED_877 ,
										MUX_10_1_IN_6 => UNWINDOWED_877 ,
										MUX_10_1_IN_7 => UNWINDOWED_1004 ,
										MUX_10_1_IN_8 => UNWINDOWED_749 ,
										MUX_10_1_IN_9 => UNWINDOWED_749 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_886
									);
MUX_REORD_UNIT_887 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_887 ,
										MUX_10_1_IN_1 => UNWINDOWED_887 ,
										MUX_10_1_IN_2 => UNWINDOWED_887 ,
										MUX_10_1_IN_3 => UNWINDOWED_894 ,
										MUX_10_1_IN_4 => UNWINDOWED_879 ,
										MUX_10_1_IN_5 => UNWINDOWED_879 ,
										MUX_10_1_IN_6 => UNWINDOWED_879 ,
										MUX_10_1_IN_7 => UNWINDOWED_1006 ,
										MUX_10_1_IN_8 => UNWINDOWED_751 ,
										MUX_10_1_IN_9 => UNWINDOWED_751 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_887
									);
MUX_REORD_UNIT_888 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_888 ,
										MUX_10_1_IN_1 => UNWINDOWED_888 ,
										MUX_10_1_IN_2 => UNWINDOWED_888 ,
										MUX_10_1_IN_3 => UNWINDOWED_881 ,
										MUX_10_1_IN_4 => UNWINDOWED_881 ,
										MUX_10_1_IN_5 => UNWINDOWED_881 ,
										MUX_10_1_IN_6 => UNWINDOWED_881 ,
										MUX_10_1_IN_7 => UNWINDOWED_1008 ,
										MUX_10_1_IN_8 => UNWINDOWED_753 ,
										MUX_10_1_IN_9 => UNWINDOWED_753 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_888
									);
MUX_REORD_UNIT_889 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_889 ,
										MUX_10_1_IN_1 => UNWINDOWED_890 ,
										MUX_10_1_IN_2 => UNWINDOWED_890 ,
										MUX_10_1_IN_3 => UNWINDOWED_883 ,
										MUX_10_1_IN_4 => UNWINDOWED_883 ,
										MUX_10_1_IN_5 => UNWINDOWED_883 ,
										MUX_10_1_IN_6 => UNWINDOWED_883 ,
										MUX_10_1_IN_7 => UNWINDOWED_1010 ,
										MUX_10_1_IN_8 => UNWINDOWED_755 ,
										MUX_10_1_IN_9 => UNWINDOWED_755 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_889
									);
MUX_REORD_UNIT_890 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_890 ,
										MUX_10_1_IN_1 => UNWINDOWED_889 ,
										MUX_10_1_IN_2 => UNWINDOWED_892 ,
										MUX_10_1_IN_3 => UNWINDOWED_885 ,
										MUX_10_1_IN_4 => UNWINDOWED_885 ,
										MUX_10_1_IN_5 => UNWINDOWED_885 ,
										MUX_10_1_IN_6 => UNWINDOWED_885 ,
										MUX_10_1_IN_7 => UNWINDOWED_1012 ,
										MUX_10_1_IN_8 => UNWINDOWED_757 ,
										MUX_10_1_IN_9 => UNWINDOWED_757 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_890
									);
MUX_REORD_UNIT_891 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_891 ,
										MUX_10_1_IN_1 => UNWINDOWED_891 ,
										MUX_10_1_IN_2 => UNWINDOWED_894 ,
										MUX_10_1_IN_3 => UNWINDOWED_887 ,
										MUX_10_1_IN_4 => UNWINDOWED_887 ,
										MUX_10_1_IN_5 => UNWINDOWED_887 ,
										MUX_10_1_IN_6 => UNWINDOWED_887 ,
										MUX_10_1_IN_7 => UNWINDOWED_1014 ,
										MUX_10_1_IN_8 => UNWINDOWED_759 ,
										MUX_10_1_IN_9 => UNWINDOWED_759 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_891
									);
MUX_REORD_UNIT_892 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_892 ,
										MUX_10_1_IN_1 => UNWINDOWED_892 ,
										MUX_10_1_IN_2 => UNWINDOWED_889 ,
										MUX_10_1_IN_3 => UNWINDOWED_889 ,
										MUX_10_1_IN_4 => UNWINDOWED_889 ,
										MUX_10_1_IN_5 => UNWINDOWED_889 ,
										MUX_10_1_IN_6 => UNWINDOWED_889 ,
										MUX_10_1_IN_7 => UNWINDOWED_1016 ,
										MUX_10_1_IN_8 => UNWINDOWED_761 ,
										MUX_10_1_IN_9 => UNWINDOWED_761 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_892
									);
MUX_REORD_UNIT_893 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_893 ,
										MUX_10_1_IN_1 => UNWINDOWED_894 ,
										MUX_10_1_IN_2 => UNWINDOWED_891 ,
										MUX_10_1_IN_3 => UNWINDOWED_891 ,
										MUX_10_1_IN_4 => UNWINDOWED_891 ,
										MUX_10_1_IN_5 => UNWINDOWED_891 ,
										MUX_10_1_IN_6 => UNWINDOWED_891 ,
										MUX_10_1_IN_7 => UNWINDOWED_1018 ,
										MUX_10_1_IN_8 => UNWINDOWED_763 ,
										MUX_10_1_IN_9 => UNWINDOWED_763 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_893
									);
MUX_REORD_UNIT_894 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_894 ,
										MUX_10_1_IN_1 => UNWINDOWED_893 ,
										MUX_10_1_IN_2 => UNWINDOWED_893 ,
										MUX_10_1_IN_3 => UNWINDOWED_893 ,
										MUX_10_1_IN_4 => UNWINDOWED_893 ,
										MUX_10_1_IN_5 => UNWINDOWED_893 ,
										MUX_10_1_IN_6 => UNWINDOWED_893 ,
										MUX_10_1_IN_7 => UNWINDOWED_1020 ,
										MUX_10_1_IN_8 => UNWINDOWED_765 ,
										MUX_10_1_IN_9 => UNWINDOWED_765 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_894
									);
MUX_REORD_UNIT_895 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_895 ,
										MUX_10_1_IN_1 => UNWINDOWED_895 ,
										MUX_10_1_IN_2 => UNWINDOWED_895 ,
										MUX_10_1_IN_3 => UNWINDOWED_895 ,
										MUX_10_1_IN_4 => UNWINDOWED_895 ,
										MUX_10_1_IN_5 => UNWINDOWED_895 ,
										MUX_10_1_IN_6 => UNWINDOWED_895 ,
										MUX_10_1_IN_7 => UNWINDOWED_1022 ,
										MUX_10_1_IN_8 => UNWINDOWED_767 ,
										MUX_10_1_IN_9 => UNWINDOWED_767 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_895
									);
MUX_REORD_UNIT_896 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_896 ,
										MUX_10_1_IN_1 => UNWINDOWED_896 ,
										MUX_10_1_IN_2 => UNWINDOWED_896 ,
										MUX_10_1_IN_3 => UNWINDOWED_896 ,
										MUX_10_1_IN_4 => UNWINDOWED_896 ,
										MUX_10_1_IN_5 => UNWINDOWED_896 ,
										MUX_10_1_IN_6 => UNWINDOWED_896 ,
										MUX_10_1_IN_7 => UNWINDOWED_769 ,
										MUX_10_1_IN_8 => UNWINDOWED_769 ,
										MUX_10_1_IN_9 => UNWINDOWED_769 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_896
									);
MUX_REORD_UNIT_897 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_897 ,
										MUX_10_1_IN_1 => UNWINDOWED_898 ,
										MUX_10_1_IN_2 => UNWINDOWED_898 ,
										MUX_10_1_IN_3 => UNWINDOWED_898 ,
										MUX_10_1_IN_4 => UNWINDOWED_898 ,
										MUX_10_1_IN_5 => UNWINDOWED_898 ,
										MUX_10_1_IN_6 => UNWINDOWED_898 ,
										MUX_10_1_IN_7 => UNWINDOWED_771 ,
										MUX_10_1_IN_8 => UNWINDOWED_771 ,
										MUX_10_1_IN_9 => UNWINDOWED_771 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_897
									);
MUX_REORD_UNIT_898 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_898 ,
										MUX_10_1_IN_1 => UNWINDOWED_897 ,
										MUX_10_1_IN_2 => UNWINDOWED_900 ,
										MUX_10_1_IN_3 => UNWINDOWED_900 ,
										MUX_10_1_IN_4 => UNWINDOWED_900 ,
										MUX_10_1_IN_5 => UNWINDOWED_900 ,
										MUX_10_1_IN_6 => UNWINDOWED_900 ,
										MUX_10_1_IN_7 => UNWINDOWED_773 ,
										MUX_10_1_IN_8 => UNWINDOWED_773 ,
										MUX_10_1_IN_9 => UNWINDOWED_773 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_898
									);
MUX_REORD_UNIT_899 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_899 ,
										MUX_10_1_IN_1 => UNWINDOWED_899 ,
										MUX_10_1_IN_2 => UNWINDOWED_902 ,
										MUX_10_1_IN_3 => UNWINDOWED_902 ,
										MUX_10_1_IN_4 => UNWINDOWED_902 ,
										MUX_10_1_IN_5 => UNWINDOWED_902 ,
										MUX_10_1_IN_6 => UNWINDOWED_902 ,
										MUX_10_1_IN_7 => UNWINDOWED_775 ,
										MUX_10_1_IN_8 => UNWINDOWED_775 ,
										MUX_10_1_IN_9 => UNWINDOWED_775 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_899
									);
MUX_REORD_UNIT_900 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_900 ,
										MUX_10_1_IN_1 => UNWINDOWED_900 ,
										MUX_10_1_IN_2 => UNWINDOWED_897 ,
										MUX_10_1_IN_3 => UNWINDOWED_904 ,
										MUX_10_1_IN_4 => UNWINDOWED_904 ,
										MUX_10_1_IN_5 => UNWINDOWED_904 ,
										MUX_10_1_IN_6 => UNWINDOWED_904 ,
										MUX_10_1_IN_7 => UNWINDOWED_777 ,
										MUX_10_1_IN_8 => UNWINDOWED_777 ,
										MUX_10_1_IN_9 => UNWINDOWED_777 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_900
									);
MUX_REORD_UNIT_901 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_901 ,
										MUX_10_1_IN_1 => UNWINDOWED_902 ,
										MUX_10_1_IN_2 => UNWINDOWED_899 ,
										MUX_10_1_IN_3 => UNWINDOWED_906 ,
										MUX_10_1_IN_4 => UNWINDOWED_906 ,
										MUX_10_1_IN_5 => UNWINDOWED_906 ,
										MUX_10_1_IN_6 => UNWINDOWED_906 ,
										MUX_10_1_IN_7 => UNWINDOWED_779 ,
										MUX_10_1_IN_8 => UNWINDOWED_779 ,
										MUX_10_1_IN_9 => UNWINDOWED_779 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_901
									);
MUX_REORD_UNIT_902 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_902 ,
										MUX_10_1_IN_1 => UNWINDOWED_901 ,
										MUX_10_1_IN_2 => UNWINDOWED_901 ,
										MUX_10_1_IN_3 => UNWINDOWED_908 ,
										MUX_10_1_IN_4 => UNWINDOWED_908 ,
										MUX_10_1_IN_5 => UNWINDOWED_908 ,
										MUX_10_1_IN_6 => UNWINDOWED_908 ,
										MUX_10_1_IN_7 => UNWINDOWED_781 ,
										MUX_10_1_IN_8 => UNWINDOWED_781 ,
										MUX_10_1_IN_9 => UNWINDOWED_781 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_902
									);
MUX_REORD_UNIT_903 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_903 ,
										MUX_10_1_IN_1 => UNWINDOWED_903 ,
										MUX_10_1_IN_2 => UNWINDOWED_903 ,
										MUX_10_1_IN_3 => UNWINDOWED_910 ,
										MUX_10_1_IN_4 => UNWINDOWED_910 ,
										MUX_10_1_IN_5 => UNWINDOWED_910 ,
										MUX_10_1_IN_6 => UNWINDOWED_910 ,
										MUX_10_1_IN_7 => UNWINDOWED_783 ,
										MUX_10_1_IN_8 => UNWINDOWED_783 ,
										MUX_10_1_IN_9 => UNWINDOWED_783 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_903
									);
MUX_REORD_UNIT_904 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_904 ,
										MUX_10_1_IN_1 => UNWINDOWED_904 ,
										MUX_10_1_IN_2 => UNWINDOWED_904 ,
										MUX_10_1_IN_3 => UNWINDOWED_897 ,
										MUX_10_1_IN_4 => UNWINDOWED_912 ,
										MUX_10_1_IN_5 => UNWINDOWED_912 ,
										MUX_10_1_IN_6 => UNWINDOWED_912 ,
										MUX_10_1_IN_7 => UNWINDOWED_785 ,
										MUX_10_1_IN_8 => UNWINDOWED_785 ,
										MUX_10_1_IN_9 => UNWINDOWED_785 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_904
									);
MUX_REORD_UNIT_905 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_905 ,
										MUX_10_1_IN_1 => UNWINDOWED_906 ,
										MUX_10_1_IN_2 => UNWINDOWED_906 ,
										MUX_10_1_IN_3 => UNWINDOWED_899 ,
										MUX_10_1_IN_4 => UNWINDOWED_914 ,
										MUX_10_1_IN_5 => UNWINDOWED_914 ,
										MUX_10_1_IN_6 => UNWINDOWED_914 ,
										MUX_10_1_IN_7 => UNWINDOWED_787 ,
										MUX_10_1_IN_8 => UNWINDOWED_787 ,
										MUX_10_1_IN_9 => UNWINDOWED_787 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_905
									);
MUX_REORD_UNIT_906 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_906 ,
										MUX_10_1_IN_1 => UNWINDOWED_905 ,
										MUX_10_1_IN_2 => UNWINDOWED_908 ,
										MUX_10_1_IN_3 => UNWINDOWED_901 ,
										MUX_10_1_IN_4 => UNWINDOWED_916 ,
										MUX_10_1_IN_5 => UNWINDOWED_916 ,
										MUX_10_1_IN_6 => UNWINDOWED_916 ,
										MUX_10_1_IN_7 => UNWINDOWED_789 ,
										MUX_10_1_IN_8 => UNWINDOWED_789 ,
										MUX_10_1_IN_9 => UNWINDOWED_789 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_906
									);
MUX_REORD_UNIT_907 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_907 ,
										MUX_10_1_IN_1 => UNWINDOWED_907 ,
										MUX_10_1_IN_2 => UNWINDOWED_910 ,
										MUX_10_1_IN_3 => UNWINDOWED_903 ,
										MUX_10_1_IN_4 => UNWINDOWED_918 ,
										MUX_10_1_IN_5 => UNWINDOWED_918 ,
										MUX_10_1_IN_6 => UNWINDOWED_918 ,
										MUX_10_1_IN_7 => UNWINDOWED_791 ,
										MUX_10_1_IN_8 => UNWINDOWED_791 ,
										MUX_10_1_IN_9 => UNWINDOWED_791 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_907
									);
MUX_REORD_UNIT_908 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_908 ,
										MUX_10_1_IN_1 => UNWINDOWED_908 ,
										MUX_10_1_IN_2 => UNWINDOWED_905 ,
										MUX_10_1_IN_3 => UNWINDOWED_905 ,
										MUX_10_1_IN_4 => UNWINDOWED_920 ,
										MUX_10_1_IN_5 => UNWINDOWED_920 ,
										MUX_10_1_IN_6 => UNWINDOWED_920 ,
										MUX_10_1_IN_7 => UNWINDOWED_793 ,
										MUX_10_1_IN_8 => UNWINDOWED_793 ,
										MUX_10_1_IN_9 => UNWINDOWED_793 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_908
									);
MUX_REORD_UNIT_909 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_909 ,
										MUX_10_1_IN_1 => UNWINDOWED_910 ,
										MUX_10_1_IN_2 => UNWINDOWED_907 ,
										MUX_10_1_IN_3 => UNWINDOWED_907 ,
										MUX_10_1_IN_4 => UNWINDOWED_922 ,
										MUX_10_1_IN_5 => UNWINDOWED_922 ,
										MUX_10_1_IN_6 => UNWINDOWED_922 ,
										MUX_10_1_IN_7 => UNWINDOWED_795 ,
										MUX_10_1_IN_8 => UNWINDOWED_795 ,
										MUX_10_1_IN_9 => UNWINDOWED_795 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_909
									);
MUX_REORD_UNIT_910 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_910 ,
										MUX_10_1_IN_1 => UNWINDOWED_909 ,
										MUX_10_1_IN_2 => UNWINDOWED_909 ,
										MUX_10_1_IN_3 => UNWINDOWED_909 ,
										MUX_10_1_IN_4 => UNWINDOWED_924 ,
										MUX_10_1_IN_5 => UNWINDOWED_924 ,
										MUX_10_1_IN_6 => UNWINDOWED_924 ,
										MUX_10_1_IN_7 => UNWINDOWED_797 ,
										MUX_10_1_IN_8 => UNWINDOWED_797 ,
										MUX_10_1_IN_9 => UNWINDOWED_797 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_910
									);
MUX_REORD_UNIT_911 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_911 ,
										MUX_10_1_IN_1 => UNWINDOWED_911 ,
										MUX_10_1_IN_2 => UNWINDOWED_911 ,
										MUX_10_1_IN_3 => UNWINDOWED_911 ,
										MUX_10_1_IN_4 => UNWINDOWED_926 ,
										MUX_10_1_IN_5 => UNWINDOWED_926 ,
										MUX_10_1_IN_6 => UNWINDOWED_926 ,
										MUX_10_1_IN_7 => UNWINDOWED_799 ,
										MUX_10_1_IN_8 => UNWINDOWED_799 ,
										MUX_10_1_IN_9 => UNWINDOWED_799 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_911
									);
MUX_REORD_UNIT_912 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_912 ,
										MUX_10_1_IN_1 => UNWINDOWED_912 ,
										MUX_10_1_IN_2 => UNWINDOWED_912 ,
										MUX_10_1_IN_3 => UNWINDOWED_912 ,
										MUX_10_1_IN_4 => UNWINDOWED_897 ,
										MUX_10_1_IN_5 => UNWINDOWED_928 ,
										MUX_10_1_IN_6 => UNWINDOWED_928 ,
										MUX_10_1_IN_7 => UNWINDOWED_801 ,
										MUX_10_1_IN_8 => UNWINDOWED_801 ,
										MUX_10_1_IN_9 => UNWINDOWED_801 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_912
									);
MUX_REORD_UNIT_913 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_913 ,
										MUX_10_1_IN_1 => UNWINDOWED_914 ,
										MUX_10_1_IN_2 => UNWINDOWED_914 ,
										MUX_10_1_IN_3 => UNWINDOWED_914 ,
										MUX_10_1_IN_4 => UNWINDOWED_899 ,
										MUX_10_1_IN_5 => UNWINDOWED_930 ,
										MUX_10_1_IN_6 => UNWINDOWED_930 ,
										MUX_10_1_IN_7 => UNWINDOWED_803 ,
										MUX_10_1_IN_8 => UNWINDOWED_803 ,
										MUX_10_1_IN_9 => UNWINDOWED_803 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_913
									);
MUX_REORD_UNIT_914 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_914 ,
										MUX_10_1_IN_1 => UNWINDOWED_913 ,
										MUX_10_1_IN_2 => UNWINDOWED_916 ,
										MUX_10_1_IN_3 => UNWINDOWED_916 ,
										MUX_10_1_IN_4 => UNWINDOWED_901 ,
										MUX_10_1_IN_5 => UNWINDOWED_932 ,
										MUX_10_1_IN_6 => UNWINDOWED_932 ,
										MUX_10_1_IN_7 => UNWINDOWED_805 ,
										MUX_10_1_IN_8 => UNWINDOWED_805 ,
										MUX_10_1_IN_9 => UNWINDOWED_805 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_914
									);
MUX_REORD_UNIT_915 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_915 ,
										MUX_10_1_IN_1 => UNWINDOWED_915 ,
										MUX_10_1_IN_2 => UNWINDOWED_918 ,
										MUX_10_1_IN_3 => UNWINDOWED_918 ,
										MUX_10_1_IN_4 => UNWINDOWED_903 ,
										MUX_10_1_IN_5 => UNWINDOWED_934 ,
										MUX_10_1_IN_6 => UNWINDOWED_934 ,
										MUX_10_1_IN_7 => UNWINDOWED_807 ,
										MUX_10_1_IN_8 => UNWINDOWED_807 ,
										MUX_10_1_IN_9 => UNWINDOWED_807 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_915
									);
MUX_REORD_UNIT_916 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_916 ,
										MUX_10_1_IN_1 => UNWINDOWED_916 ,
										MUX_10_1_IN_2 => UNWINDOWED_913 ,
										MUX_10_1_IN_3 => UNWINDOWED_920 ,
										MUX_10_1_IN_4 => UNWINDOWED_905 ,
										MUX_10_1_IN_5 => UNWINDOWED_936 ,
										MUX_10_1_IN_6 => UNWINDOWED_936 ,
										MUX_10_1_IN_7 => UNWINDOWED_809 ,
										MUX_10_1_IN_8 => UNWINDOWED_809 ,
										MUX_10_1_IN_9 => UNWINDOWED_809 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_916
									);
MUX_REORD_UNIT_917 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_917 ,
										MUX_10_1_IN_1 => UNWINDOWED_918 ,
										MUX_10_1_IN_2 => UNWINDOWED_915 ,
										MUX_10_1_IN_3 => UNWINDOWED_922 ,
										MUX_10_1_IN_4 => UNWINDOWED_907 ,
										MUX_10_1_IN_5 => UNWINDOWED_938 ,
										MUX_10_1_IN_6 => UNWINDOWED_938 ,
										MUX_10_1_IN_7 => UNWINDOWED_811 ,
										MUX_10_1_IN_8 => UNWINDOWED_811 ,
										MUX_10_1_IN_9 => UNWINDOWED_811 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_917
									);
MUX_REORD_UNIT_918 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_918 ,
										MUX_10_1_IN_1 => UNWINDOWED_917 ,
										MUX_10_1_IN_2 => UNWINDOWED_917 ,
										MUX_10_1_IN_3 => UNWINDOWED_924 ,
										MUX_10_1_IN_4 => UNWINDOWED_909 ,
										MUX_10_1_IN_5 => UNWINDOWED_940 ,
										MUX_10_1_IN_6 => UNWINDOWED_940 ,
										MUX_10_1_IN_7 => UNWINDOWED_813 ,
										MUX_10_1_IN_8 => UNWINDOWED_813 ,
										MUX_10_1_IN_9 => UNWINDOWED_813 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_918
									);
MUX_REORD_UNIT_919 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_919 ,
										MUX_10_1_IN_1 => UNWINDOWED_919 ,
										MUX_10_1_IN_2 => UNWINDOWED_919 ,
										MUX_10_1_IN_3 => UNWINDOWED_926 ,
										MUX_10_1_IN_4 => UNWINDOWED_911 ,
										MUX_10_1_IN_5 => UNWINDOWED_942 ,
										MUX_10_1_IN_6 => UNWINDOWED_942 ,
										MUX_10_1_IN_7 => UNWINDOWED_815 ,
										MUX_10_1_IN_8 => UNWINDOWED_815 ,
										MUX_10_1_IN_9 => UNWINDOWED_815 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_919
									);
MUX_REORD_UNIT_920 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_920 ,
										MUX_10_1_IN_1 => UNWINDOWED_920 ,
										MUX_10_1_IN_2 => UNWINDOWED_920 ,
										MUX_10_1_IN_3 => UNWINDOWED_913 ,
										MUX_10_1_IN_4 => UNWINDOWED_913 ,
										MUX_10_1_IN_5 => UNWINDOWED_944 ,
										MUX_10_1_IN_6 => UNWINDOWED_944 ,
										MUX_10_1_IN_7 => UNWINDOWED_817 ,
										MUX_10_1_IN_8 => UNWINDOWED_817 ,
										MUX_10_1_IN_9 => UNWINDOWED_817 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_920
									);
MUX_REORD_UNIT_921 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_921 ,
										MUX_10_1_IN_1 => UNWINDOWED_922 ,
										MUX_10_1_IN_2 => UNWINDOWED_922 ,
										MUX_10_1_IN_3 => UNWINDOWED_915 ,
										MUX_10_1_IN_4 => UNWINDOWED_915 ,
										MUX_10_1_IN_5 => UNWINDOWED_946 ,
										MUX_10_1_IN_6 => UNWINDOWED_946 ,
										MUX_10_1_IN_7 => UNWINDOWED_819 ,
										MUX_10_1_IN_8 => UNWINDOWED_819 ,
										MUX_10_1_IN_9 => UNWINDOWED_819 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_921
									);
MUX_REORD_UNIT_922 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_922 ,
										MUX_10_1_IN_1 => UNWINDOWED_921 ,
										MUX_10_1_IN_2 => UNWINDOWED_924 ,
										MUX_10_1_IN_3 => UNWINDOWED_917 ,
										MUX_10_1_IN_4 => UNWINDOWED_917 ,
										MUX_10_1_IN_5 => UNWINDOWED_948 ,
										MUX_10_1_IN_6 => UNWINDOWED_948 ,
										MUX_10_1_IN_7 => UNWINDOWED_821 ,
										MUX_10_1_IN_8 => UNWINDOWED_821 ,
										MUX_10_1_IN_9 => UNWINDOWED_821 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_922
									);
MUX_REORD_UNIT_923 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_923 ,
										MUX_10_1_IN_1 => UNWINDOWED_923 ,
										MUX_10_1_IN_2 => UNWINDOWED_926 ,
										MUX_10_1_IN_3 => UNWINDOWED_919 ,
										MUX_10_1_IN_4 => UNWINDOWED_919 ,
										MUX_10_1_IN_5 => UNWINDOWED_950 ,
										MUX_10_1_IN_6 => UNWINDOWED_950 ,
										MUX_10_1_IN_7 => UNWINDOWED_823 ,
										MUX_10_1_IN_8 => UNWINDOWED_823 ,
										MUX_10_1_IN_9 => UNWINDOWED_823 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_923
									);
MUX_REORD_UNIT_924 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_924 ,
										MUX_10_1_IN_1 => UNWINDOWED_924 ,
										MUX_10_1_IN_2 => UNWINDOWED_921 ,
										MUX_10_1_IN_3 => UNWINDOWED_921 ,
										MUX_10_1_IN_4 => UNWINDOWED_921 ,
										MUX_10_1_IN_5 => UNWINDOWED_952 ,
										MUX_10_1_IN_6 => UNWINDOWED_952 ,
										MUX_10_1_IN_7 => UNWINDOWED_825 ,
										MUX_10_1_IN_8 => UNWINDOWED_825 ,
										MUX_10_1_IN_9 => UNWINDOWED_825 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_924
									);
MUX_REORD_UNIT_925 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_925 ,
										MUX_10_1_IN_1 => UNWINDOWED_926 ,
										MUX_10_1_IN_2 => UNWINDOWED_923 ,
										MUX_10_1_IN_3 => UNWINDOWED_923 ,
										MUX_10_1_IN_4 => UNWINDOWED_923 ,
										MUX_10_1_IN_5 => UNWINDOWED_954 ,
										MUX_10_1_IN_6 => UNWINDOWED_954 ,
										MUX_10_1_IN_7 => UNWINDOWED_827 ,
										MUX_10_1_IN_8 => UNWINDOWED_827 ,
										MUX_10_1_IN_9 => UNWINDOWED_827 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_925
									);
MUX_REORD_UNIT_926 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_926 ,
										MUX_10_1_IN_1 => UNWINDOWED_925 ,
										MUX_10_1_IN_2 => UNWINDOWED_925 ,
										MUX_10_1_IN_3 => UNWINDOWED_925 ,
										MUX_10_1_IN_4 => UNWINDOWED_925 ,
										MUX_10_1_IN_5 => UNWINDOWED_956 ,
										MUX_10_1_IN_6 => UNWINDOWED_956 ,
										MUX_10_1_IN_7 => UNWINDOWED_829 ,
										MUX_10_1_IN_8 => UNWINDOWED_829 ,
										MUX_10_1_IN_9 => UNWINDOWED_829 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_926
									);
MUX_REORD_UNIT_927 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_927 ,
										MUX_10_1_IN_1 => UNWINDOWED_927 ,
										MUX_10_1_IN_2 => UNWINDOWED_927 ,
										MUX_10_1_IN_3 => UNWINDOWED_927 ,
										MUX_10_1_IN_4 => UNWINDOWED_927 ,
										MUX_10_1_IN_5 => UNWINDOWED_958 ,
										MUX_10_1_IN_6 => UNWINDOWED_958 ,
										MUX_10_1_IN_7 => UNWINDOWED_831 ,
										MUX_10_1_IN_8 => UNWINDOWED_831 ,
										MUX_10_1_IN_9 => UNWINDOWED_831 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_927
									);
MUX_REORD_UNIT_928 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_928 ,
										MUX_10_1_IN_1 => UNWINDOWED_928 ,
										MUX_10_1_IN_2 => UNWINDOWED_928 ,
										MUX_10_1_IN_3 => UNWINDOWED_928 ,
										MUX_10_1_IN_4 => UNWINDOWED_928 ,
										MUX_10_1_IN_5 => UNWINDOWED_897 ,
										MUX_10_1_IN_6 => UNWINDOWED_960 ,
										MUX_10_1_IN_7 => UNWINDOWED_833 ,
										MUX_10_1_IN_8 => UNWINDOWED_833 ,
										MUX_10_1_IN_9 => UNWINDOWED_833 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_928
									);
MUX_REORD_UNIT_929 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_929 ,
										MUX_10_1_IN_1 => UNWINDOWED_930 ,
										MUX_10_1_IN_2 => UNWINDOWED_930 ,
										MUX_10_1_IN_3 => UNWINDOWED_930 ,
										MUX_10_1_IN_4 => UNWINDOWED_930 ,
										MUX_10_1_IN_5 => UNWINDOWED_899 ,
										MUX_10_1_IN_6 => UNWINDOWED_962 ,
										MUX_10_1_IN_7 => UNWINDOWED_835 ,
										MUX_10_1_IN_8 => UNWINDOWED_835 ,
										MUX_10_1_IN_9 => UNWINDOWED_835 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_929
									);
MUX_REORD_UNIT_930 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_930 ,
										MUX_10_1_IN_1 => UNWINDOWED_929 ,
										MUX_10_1_IN_2 => UNWINDOWED_932 ,
										MUX_10_1_IN_3 => UNWINDOWED_932 ,
										MUX_10_1_IN_4 => UNWINDOWED_932 ,
										MUX_10_1_IN_5 => UNWINDOWED_901 ,
										MUX_10_1_IN_6 => UNWINDOWED_964 ,
										MUX_10_1_IN_7 => UNWINDOWED_837 ,
										MUX_10_1_IN_8 => UNWINDOWED_837 ,
										MUX_10_1_IN_9 => UNWINDOWED_837 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_930
									);
MUX_REORD_UNIT_931 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_931 ,
										MUX_10_1_IN_1 => UNWINDOWED_931 ,
										MUX_10_1_IN_2 => UNWINDOWED_934 ,
										MUX_10_1_IN_3 => UNWINDOWED_934 ,
										MUX_10_1_IN_4 => UNWINDOWED_934 ,
										MUX_10_1_IN_5 => UNWINDOWED_903 ,
										MUX_10_1_IN_6 => UNWINDOWED_966 ,
										MUX_10_1_IN_7 => UNWINDOWED_839 ,
										MUX_10_1_IN_8 => UNWINDOWED_839 ,
										MUX_10_1_IN_9 => UNWINDOWED_839 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_931
									);
MUX_REORD_UNIT_932 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_932 ,
										MUX_10_1_IN_1 => UNWINDOWED_932 ,
										MUX_10_1_IN_2 => UNWINDOWED_929 ,
										MUX_10_1_IN_3 => UNWINDOWED_936 ,
										MUX_10_1_IN_4 => UNWINDOWED_936 ,
										MUX_10_1_IN_5 => UNWINDOWED_905 ,
										MUX_10_1_IN_6 => UNWINDOWED_968 ,
										MUX_10_1_IN_7 => UNWINDOWED_841 ,
										MUX_10_1_IN_8 => UNWINDOWED_841 ,
										MUX_10_1_IN_9 => UNWINDOWED_841 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_932
									);
MUX_REORD_UNIT_933 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_933 ,
										MUX_10_1_IN_1 => UNWINDOWED_934 ,
										MUX_10_1_IN_2 => UNWINDOWED_931 ,
										MUX_10_1_IN_3 => UNWINDOWED_938 ,
										MUX_10_1_IN_4 => UNWINDOWED_938 ,
										MUX_10_1_IN_5 => UNWINDOWED_907 ,
										MUX_10_1_IN_6 => UNWINDOWED_970 ,
										MUX_10_1_IN_7 => UNWINDOWED_843 ,
										MUX_10_1_IN_8 => UNWINDOWED_843 ,
										MUX_10_1_IN_9 => UNWINDOWED_843 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_933
									);
MUX_REORD_UNIT_934 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_934 ,
										MUX_10_1_IN_1 => UNWINDOWED_933 ,
										MUX_10_1_IN_2 => UNWINDOWED_933 ,
										MUX_10_1_IN_3 => UNWINDOWED_940 ,
										MUX_10_1_IN_4 => UNWINDOWED_940 ,
										MUX_10_1_IN_5 => UNWINDOWED_909 ,
										MUX_10_1_IN_6 => UNWINDOWED_972 ,
										MUX_10_1_IN_7 => UNWINDOWED_845 ,
										MUX_10_1_IN_8 => UNWINDOWED_845 ,
										MUX_10_1_IN_9 => UNWINDOWED_845 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_934
									);
MUX_REORD_UNIT_935 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_935 ,
										MUX_10_1_IN_1 => UNWINDOWED_935 ,
										MUX_10_1_IN_2 => UNWINDOWED_935 ,
										MUX_10_1_IN_3 => UNWINDOWED_942 ,
										MUX_10_1_IN_4 => UNWINDOWED_942 ,
										MUX_10_1_IN_5 => UNWINDOWED_911 ,
										MUX_10_1_IN_6 => UNWINDOWED_974 ,
										MUX_10_1_IN_7 => UNWINDOWED_847 ,
										MUX_10_1_IN_8 => UNWINDOWED_847 ,
										MUX_10_1_IN_9 => UNWINDOWED_847 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_935
									);
MUX_REORD_UNIT_936 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_936 ,
										MUX_10_1_IN_1 => UNWINDOWED_936 ,
										MUX_10_1_IN_2 => UNWINDOWED_936 ,
										MUX_10_1_IN_3 => UNWINDOWED_929 ,
										MUX_10_1_IN_4 => UNWINDOWED_944 ,
										MUX_10_1_IN_5 => UNWINDOWED_913 ,
										MUX_10_1_IN_6 => UNWINDOWED_976 ,
										MUX_10_1_IN_7 => UNWINDOWED_849 ,
										MUX_10_1_IN_8 => UNWINDOWED_849 ,
										MUX_10_1_IN_9 => UNWINDOWED_849 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_936
									);
MUX_REORD_UNIT_937 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_937 ,
										MUX_10_1_IN_1 => UNWINDOWED_938 ,
										MUX_10_1_IN_2 => UNWINDOWED_938 ,
										MUX_10_1_IN_3 => UNWINDOWED_931 ,
										MUX_10_1_IN_4 => UNWINDOWED_946 ,
										MUX_10_1_IN_5 => UNWINDOWED_915 ,
										MUX_10_1_IN_6 => UNWINDOWED_978 ,
										MUX_10_1_IN_7 => UNWINDOWED_851 ,
										MUX_10_1_IN_8 => UNWINDOWED_851 ,
										MUX_10_1_IN_9 => UNWINDOWED_851 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_937
									);
MUX_REORD_UNIT_938 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_938 ,
										MUX_10_1_IN_1 => UNWINDOWED_937 ,
										MUX_10_1_IN_2 => UNWINDOWED_940 ,
										MUX_10_1_IN_3 => UNWINDOWED_933 ,
										MUX_10_1_IN_4 => UNWINDOWED_948 ,
										MUX_10_1_IN_5 => UNWINDOWED_917 ,
										MUX_10_1_IN_6 => UNWINDOWED_980 ,
										MUX_10_1_IN_7 => UNWINDOWED_853 ,
										MUX_10_1_IN_8 => UNWINDOWED_853 ,
										MUX_10_1_IN_9 => UNWINDOWED_853 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_938
									);
MUX_REORD_UNIT_939 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_939 ,
										MUX_10_1_IN_1 => UNWINDOWED_939 ,
										MUX_10_1_IN_2 => UNWINDOWED_942 ,
										MUX_10_1_IN_3 => UNWINDOWED_935 ,
										MUX_10_1_IN_4 => UNWINDOWED_950 ,
										MUX_10_1_IN_5 => UNWINDOWED_919 ,
										MUX_10_1_IN_6 => UNWINDOWED_982 ,
										MUX_10_1_IN_7 => UNWINDOWED_855 ,
										MUX_10_1_IN_8 => UNWINDOWED_855 ,
										MUX_10_1_IN_9 => UNWINDOWED_855 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_939
									);
MUX_REORD_UNIT_940 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_940 ,
										MUX_10_1_IN_1 => UNWINDOWED_940 ,
										MUX_10_1_IN_2 => UNWINDOWED_937 ,
										MUX_10_1_IN_3 => UNWINDOWED_937 ,
										MUX_10_1_IN_4 => UNWINDOWED_952 ,
										MUX_10_1_IN_5 => UNWINDOWED_921 ,
										MUX_10_1_IN_6 => UNWINDOWED_984 ,
										MUX_10_1_IN_7 => UNWINDOWED_857 ,
										MUX_10_1_IN_8 => UNWINDOWED_857 ,
										MUX_10_1_IN_9 => UNWINDOWED_857 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_940
									);
MUX_REORD_UNIT_941 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_941 ,
										MUX_10_1_IN_1 => UNWINDOWED_942 ,
										MUX_10_1_IN_2 => UNWINDOWED_939 ,
										MUX_10_1_IN_3 => UNWINDOWED_939 ,
										MUX_10_1_IN_4 => UNWINDOWED_954 ,
										MUX_10_1_IN_5 => UNWINDOWED_923 ,
										MUX_10_1_IN_6 => UNWINDOWED_986 ,
										MUX_10_1_IN_7 => UNWINDOWED_859 ,
										MUX_10_1_IN_8 => UNWINDOWED_859 ,
										MUX_10_1_IN_9 => UNWINDOWED_859 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_941
									);
MUX_REORD_UNIT_942 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_942 ,
										MUX_10_1_IN_1 => UNWINDOWED_941 ,
										MUX_10_1_IN_2 => UNWINDOWED_941 ,
										MUX_10_1_IN_3 => UNWINDOWED_941 ,
										MUX_10_1_IN_4 => UNWINDOWED_956 ,
										MUX_10_1_IN_5 => UNWINDOWED_925 ,
										MUX_10_1_IN_6 => UNWINDOWED_988 ,
										MUX_10_1_IN_7 => UNWINDOWED_861 ,
										MUX_10_1_IN_8 => UNWINDOWED_861 ,
										MUX_10_1_IN_9 => UNWINDOWED_861 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_942
									);
MUX_REORD_UNIT_943 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_943 ,
										MUX_10_1_IN_1 => UNWINDOWED_943 ,
										MUX_10_1_IN_2 => UNWINDOWED_943 ,
										MUX_10_1_IN_3 => UNWINDOWED_943 ,
										MUX_10_1_IN_4 => UNWINDOWED_958 ,
										MUX_10_1_IN_5 => UNWINDOWED_927 ,
										MUX_10_1_IN_6 => UNWINDOWED_990 ,
										MUX_10_1_IN_7 => UNWINDOWED_863 ,
										MUX_10_1_IN_8 => UNWINDOWED_863 ,
										MUX_10_1_IN_9 => UNWINDOWED_863 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_943
									);
MUX_REORD_UNIT_944 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_944 ,
										MUX_10_1_IN_1 => UNWINDOWED_944 ,
										MUX_10_1_IN_2 => UNWINDOWED_944 ,
										MUX_10_1_IN_3 => UNWINDOWED_944 ,
										MUX_10_1_IN_4 => UNWINDOWED_929 ,
										MUX_10_1_IN_5 => UNWINDOWED_929 ,
										MUX_10_1_IN_6 => UNWINDOWED_992 ,
										MUX_10_1_IN_7 => UNWINDOWED_865 ,
										MUX_10_1_IN_8 => UNWINDOWED_865 ,
										MUX_10_1_IN_9 => UNWINDOWED_865 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_944
									);
MUX_REORD_UNIT_945 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_945 ,
										MUX_10_1_IN_1 => UNWINDOWED_946 ,
										MUX_10_1_IN_2 => UNWINDOWED_946 ,
										MUX_10_1_IN_3 => UNWINDOWED_946 ,
										MUX_10_1_IN_4 => UNWINDOWED_931 ,
										MUX_10_1_IN_5 => UNWINDOWED_931 ,
										MUX_10_1_IN_6 => UNWINDOWED_994 ,
										MUX_10_1_IN_7 => UNWINDOWED_867 ,
										MUX_10_1_IN_8 => UNWINDOWED_867 ,
										MUX_10_1_IN_9 => UNWINDOWED_867 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_945
									);
MUX_REORD_UNIT_946 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_946 ,
										MUX_10_1_IN_1 => UNWINDOWED_945 ,
										MUX_10_1_IN_2 => UNWINDOWED_948 ,
										MUX_10_1_IN_3 => UNWINDOWED_948 ,
										MUX_10_1_IN_4 => UNWINDOWED_933 ,
										MUX_10_1_IN_5 => UNWINDOWED_933 ,
										MUX_10_1_IN_6 => UNWINDOWED_996 ,
										MUX_10_1_IN_7 => UNWINDOWED_869 ,
										MUX_10_1_IN_8 => UNWINDOWED_869 ,
										MUX_10_1_IN_9 => UNWINDOWED_869 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_946
									);
MUX_REORD_UNIT_947 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_947 ,
										MUX_10_1_IN_1 => UNWINDOWED_947 ,
										MUX_10_1_IN_2 => UNWINDOWED_950 ,
										MUX_10_1_IN_3 => UNWINDOWED_950 ,
										MUX_10_1_IN_4 => UNWINDOWED_935 ,
										MUX_10_1_IN_5 => UNWINDOWED_935 ,
										MUX_10_1_IN_6 => UNWINDOWED_998 ,
										MUX_10_1_IN_7 => UNWINDOWED_871 ,
										MUX_10_1_IN_8 => UNWINDOWED_871 ,
										MUX_10_1_IN_9 => UNWINDOWED_871 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_947
									);
MUX_REORD_UNIT_948 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_948 ,
										MUX_10_1_IN_1 => UNWINDOWED_948 ,
										MUX_10_1_IN_2 => UNWINDOWED_945 ,
										MUX_10_1_IN_3 => UNWINDOWED_952 ,
										MUX_10_1_IN_4 => UNWINDOWED_937 ,
										MUX_10_1_IN_5 => UNWINDOWED_937 ,
										MUX_10_1_IN_6 => UNWINDOWED_1000 ,
										MUX_10_1_IN_7 => UNWINDOWED_873 ,
										MUX_10_1_IN_8 => UNWINDOWED_873 ,
										MUX_10_1_IN_9 => UNWINDOWED_873 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_948
									);
MUX_REORD_UNIT_949 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_949 ,
										MUX_10_1_IN_1 => UNWINDOWED_950 ,
										MUX_10_1_IN_2 => UNWINDOWED_947 ,
										MUX_10_1_IN_3 => UNWINDOWED_954 ,
										MUX_10_1_IN_4 => UNWINDOWED_939 ,
										MUX_10_1_IN_5 => UNWINDOWED_939 ,
										MUX_10_1_IN_6 => UNWINDOWED_1002 ,
										MUX_10_1_IN_7 => UNWINDOWED_875 ,
										MUX_10_1_IN_8 => UNWINDOWED_875 ,
										MUX_10_1_IN_9 => UNWINDOWED_875 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_949
									);
MUX_REORD_UNIT_950 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_950 ,
										MUX_10_1_IN_1 => UNWINDOWED_949 ,
										MUX_10_1_IN_2 => UNWINDOWED_949 ,
										MUX_10_1_IN_3 => UNWINDOWED_956 ,
										MUX_10_1_IN_4 => UNWINDOWED_941 ,
										MUX_10_1_IN_5 => UNWINDOWED_941 ,
										MUX_10_1_IN_6 => UNWINDOWED_1004 ,
										MUX_10_1_IN_7 => UNWINDOWED_877 ,
										MUX_10_1_IN_8 => UNWINDOWED_877 ,
										MUX_10_1_IN_9 => UNWINDOWED_877 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_950
									);
MUX_REORD_UNIT_951 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_951 ,
										MUX_10_1_IN_1 => UNWINDOWED_951 ,
										MUX_10_1_IN_2 => UNWINDOWED_951 ,
										MUX_10_1_IN_3 => UNWINDOWED_958 ,
										MUX_10_1_IN_4 => UNWINDOWED_943 ,
										MUX_10_1_IN_5 => UNWINDOWED_943 ,
										MUX_10_1_IN_6 => UNWINDOWED_1006 ,
										MUX_10_1_IN_7 => UNWINDOWED_879 ,
										MUX_10_1_IN_8 => UNWINDOWED_879 ,
										MUX_10_1_IN_9 => UNWINDOWED_879 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_951
									);
MUX_REORD_UNIT_952 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_952 ,
										MUX_10_1_IN_1 => UNWINDOWED_952 ,
										MUX_10_1_IN_2 => UNWINDOWED_952 ,
										MUX_10_1_IN_3 => UNWINDOWED_945 ,
										MUX_10_1_IN_4 => UNWINDOWED_945 ,
										MUX_10_1_IN_5 => UNWINDOWED_945 ,
										MUX_10_1_IN_6 => UNWINDOWED_1008 ,
										MUX_10_1_IN_7 => UNWINDOWED_881 ,
										MUX_10_1_IN_8 => UNWINDOWED_881 ,
										MUX_10_1_IN_9 => UNWINDOWED_881 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_952
									);
MUX_REORD_UNIT_953 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_953 ,
										MUX_10_1_IN_1 => UNWINDOWED_954 ,
										MUX_10_1_IN_2 => UNWINDOWED_954 ,
										MUX_10_1_IN_3 => UNWINDOWED_947 ,
										MUX_10_1_IN_4 => UNWINDOWED_947 ,
										MUX_10_1_IN_5 => UNWINDOWED_947 ,
										MUX_10_1_IN_6 => UNWINDOWED_1010 ,
										MUX_10_1_IN_7 => UNWINDOWED_883 ,
										MUX_10_1_IN_8 => UNWINDOWED_883 ,
										MUX_10_1_IN_9 => UNWINDOWED_883 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_953
									);
MUX_REORD_UNIT_954 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_954 ,
										MUX_10_1_IN_1 => UNWINDOWED_953 ,
										MUX_10_1_IN_2 => UNWINDOWED_956 ,
										MUX_10_1_IN_3 => UNWINDOWED_949 ,
										MUX_10_1_IN_4 => UNWINDOWED_949 ,
										MUX_10_1_IN_5 => UNWINDOWED_949 ,
										MUX_10_1_IN_6 => UNWINDOWED_1012 ,
										MUX_10_1_IN_7 => UNWINDOWED_885 ,
										MUX_10_1_IN_8 => UNWINDOWED_885 ,
										MUX_10_1_IN_9 => UNWINDOWED_885 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_954
									);
MUX_REORD_UNIT_955 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_955 ,
										MUX_10_1_IN_1 => UNWINDOWED_955 ,
										MUX_10_1_IN_2 => UNWINDOWED_958 ,
										MUX_10_1_IN_3 => UNWINDOWED_951 ,
										MUX_10_1_IN_4 => UNWINDOWED_951 ,
										MUX_10_1_IN_5 => UNWINDOWED_951 ,
										MUX_10_1_IN_6 => UNWINDOWED_1014 ,
										MUX_10_1_IN_7 => UNWINDOWED_887 ,
										MUX_10_1_IN_8 => UNWINDOWED_887 ,
										MUX_10_1_IN_9 => UNWINDOWED_887 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_955
									);
MUX_REORD_UNIT_956 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_956 ,
										MUX_10_1_IN_1 => UNWINDOWED_956 ,
										MUX_10_1_IN_2 => UNWINDOWED_953 ,
										MUX_10_1_IN_3 => UNWINDOWED_953 ,
										MUX_10_1_IN_4 => UNWINDOWED_953 ,
										MUX_10_1_IN_5 => UNWINDOWED_953 ,
										MUX_10_1_IN_6 => UNWINDOWED_1016 ,
										MUX_10_1_IN_7 => UNWINDOWED_889 ,
										MUX_10_1_IN_8 => UNWINDOWED_889 ,
										MUX_10_1_IN_9 => UNWINDOWED_889 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_956
									);
MUX_REORD_UNIT_957 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_957 ,
										MUX_10_1_IN_1 => UNWINDOWED_958 ,
										MUX_10_1_IN_2 => UNWINDOWED_955 ,
										MUX_10_1_IN_3 => UNWINDOWED_955 ,
										MUX_10_1_IN_4 => UNWINDOWED_955 ,
										MUX_10_1_IN_5 => UNWINDOWED_955 ,
										MUX_10_1_IN_6 => UNWINDOWED_1018 ,
										MUX_10_1_IN_7 => UNWINDOWED_891 ,
										MUX_10_1_IN_8 => UNWINDOWED_891 ,
										MUX_10_1_IN_9 => UNWINDOWED_891 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_957
									);
MUX_REORD_UNIT_958 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_958 ,
										MUX_10_1_IN_1 => UNWINDOWED_957 ,
										MUX_10_1_IN_2 => UNWINDOWED_957 ,
										MUX_10_1_IN_3 => UNWINDOWED_957 ,
										MUX_10_1_IN_4 => UNWINDOWED_957 ,
										MUX_10_1_IN_5 => UNWINDOWED_957 ,
										MUX_10_1_IN_6 => UNWINDOWED_1020 ,
										MUX_10_1_IN_7 => UNWINDOWED_893 ,
										MUX_10_1_IN_8 => UNWINDOWED_893 ,
										MUX_10_1_IN_9 => UNWINDOWED_893 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_958
									);
MUX_REORD_UNIT_959 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_959 ,
										MUX_10_1_IN_1 => UNWINDOWED_959 ,
										MUX_10_1_IN_2 => UNWINDOWED_959 ,
										MUX_10_1_IN_3 => UNWINDOWED_959 ,
										MUX_10_1_IN_4 => UNWINDOWED_959 ,
										MUX_10_1_IN_5 => UNWINDOWED_959 ,
										MUX_10_1_IN_6 => UNWINDOWED_1022 ,
										MUX_10_1_IN_7 => UNWINDOWED_895 ,
										MUX_10_1_IN_8 => UNWINDOWED_895 ,
										MUX_10_1_IN_9 => UNWINDOWED_895 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_959
									);
MUX_REORD_UNIT_960 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_960 ,
										MUX_10_1_IN_1 => UNWINDOWED_960 ,
										MUX_10_1_IN_2 => UNWINDOWED_960 ,
										MUX_10_1_IN_3 => UNWINDOWED_960 ,
										MUX_10_1_IN_4 => UNWINDOWED_960 ,
										MUX_10_1_IN_5 => UNWINDOWED_960 ,
										MUX_10_1_IN_6 => UNWINDOWED_897 ,
										MUX_10_1_IN_7 => UNWINDOWED_897 ,
										MUX_10_1_IN_8 => UNWINDOWED_897 ,
										MUX_10_1_IN_9 => UNWINDOWED_897 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_960
									);
MUX_REORD_UNIT_961 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_961 ,
										MUX_10_1_IN_1 => UNWINDOWED_962 ,
										MUX_10_1_IN_2 => UNWINDOWED_962 ,
										MUX_10_1_IN_3 => UNWINDOWED_962 ,
										MUX_10_1_IN_4 => UNWINDOWED_962 ,
										MUX_10_1_IN_5 => UNWINDOWED_962 ,
										MUX_10_1_IN_6 => UNWINDOWED_899 ,
										MUX_10_1_IN_7 => UNWINDOWED_899 ,
										MUX_10_1_IN_8 => UNWINDOWED_899 ,
										MUX_10_1_IN_9 => UNWINDOWED_899 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_961
									);
MUX_REORD_UNIT_962 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_962 ,
										MUX_10_1_IN_1 => UNWINDOWED_961 ,
										MUX_10_1_IN_2 => UNWINDOWED_964 ,
										MUX_10_1_IN_3 => UNWINDOWED_964 ,
										MUX_10_1_IN_4 => UNWINDOWED_964 ,
										MUX_10_1_IN_5 => UNWINDOWED_964 ,
										MUX_10_1_IN_6 => UNWINDOWED_901 ,
										MUX_10_1_IN_7 => UNWINDOWED_901 ,
										MUX_10_1_IN_8 => UNWINDOWED_901 ,
										MUX_10_1_IN_9 => UNWINDOWED_901 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_962
									);
MUX_REORD_UNIT_963 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_963 ,
										MUX_10_1_IN_1 => UNWINDOWED_963 ,
										MUX_10_1_IN_2 => UNWINDOWED_966 ,
										MUX_10_1_IN_3 => UNWINDOWED_966 ,
										MUX_10_1_IN_4 => UNWINDOWED_966 ,
										MUX_10_1_IN_5 => UNWINDOWED_966 ,
										MUX_10_1_IN_6 => UNWINDOWED_903 ,
										MUX_10_1_IN_7 => UNWINDOWED_903 ,
										MUX_10_1_IN_8 => UNWINDOWED_903 ,
										MUX_10_1_IN_9 => UNWINDOWED_903 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_963
									);
MUX_REORD_UNIT_964 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_964 ,
										MUX_10_1_IN_1 => UNWINDOWED_964 ,
										MUX_10_1_IN_2 => UNWINDOWED_961 ,
										MUX_10_1_IN_3 => UNWINDOWED_968 ,
										MUX_10_1_IN_4 => UNWINDOWED_968 ,
										MUX_10_1_IN_5 => UNWINDOWED_968 ,
										MUX_10_1_IN_6 => UNWINDOWED_905 ,
										MUX_10_1_IN_7 => UNWINDOWED_905 ,
										MUX_10_1_IN_8 => UNWINDOWED_905 ,
										MUX_10_1_IN_9 => UNWINDOWED_905 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_964
									);
MUX_REORD_UNIT_965 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_965 ,
										MUX_10_1_IN_1 => UNWINDOWED_966 ,
										MUX_10_1_IN_2 => UNWINDOWED_963 ,
										MUX_10_1_IN_3 => UNWINDOWED_970 ,
										MUX_10_1_IN_4 => UNWINDOWED_970 ,
										MUX_10_1_IN_5 => UNWINDOWED_970 ,
										MUX_10_1_IN_6 => UNWINDOWED_907 ,
										MUX_10_1_IN_7 => UNWINDOWED_907 ,
										MUX_10_1_IN_8 => UNWINDOWED_907 ,
										MUX_10_1_IN_9 => UNWINDOWED_907 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_965
									);
MUX_REORD_UNIT_966 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_966 ,
										MUX_10_1_IN_1 => UNWINDOWED_965 ,
										MUX_10_1_IN_2 => UNWINDOWED_965 ,
										MUX_10_1_IN_3 => UNWINDOWED_972 ,
										MUX_10_1_IN_4 => UNWINDOWED_972 ,
										MUX_10_1_IN_5 => UNWINDOWED_972 ,
										MUX_10_1_IN_6 => UNWINDOWED_909 ,
										MUX_10_1_IN_7 => UNWINDOWED_909 ,
										MUX_10_1_IN_8 => UNWINDOWED_909 ,
										MUX_10_1_IN_9 => UNWINDOWED_909 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_966
									);
MUX_REORD_UNIT_967 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_967 ,
										MUX_10_1_IN_1 => UNWINDOWED_967 ,
										MUX_10_1_IN_2 => UNWINDOWED_967 ,
										MUX_10_1_IN_3 => UNWINDOWED_974 ,
										MUX_10_1_IN_4 => UNWINDOWED_974 ,
										MUX_10_1_IN_5 => UNWINDOWED_974 ,
										MUX_10_1_IN_6 => UNWINDOWED_911 ,
										MUX_10_1_IN_7 => UNWINDOWED_911 ,
										MUX_10_1_IN_8 => UNWINDOWED_911 ,
										MUX_10_1_IN_9 => UNWINDOWED_911 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_967
									);
MUX_REORD_UNIT_968 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_968 ,
										MUX_10_1_IN_1 => UNWINDOWED_968 ,
										MUX_10_1_IN_2 => UNWINDOWED_968 ,
										MUX_10_1_IN_3 => UNWINDOWED_961 ,
										MUX_10_1_IN_4 => UNWINDOWED_976 ,
										MUX_10_1_IN_5 => UNWINDOWED_976 ,
										MUX_10_1_IN_6 => UNWINDOWED_913 ,
										MUX_10_1_IN_7 => UNWINDOWED_913 ,
										MUX_10_1_IN_8 => UNWINDOWED_913 ,
										MUX_10_1_IN_9 => UNWINDOWED_913 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_968
									);
MUX_REORD_UNIT_969 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_969 ,
										MUX_10_1_IN_1 => UNWINDOWED_970 ,
										MUX_10_1_IN_2 => UNWINDOWED_970 ,
										MUX_10_1_IN_3 => UNWINDOWED_963 ,
										MUX_10_1_IN_4 => UNWINDOWED_978 ,
										MUX_10_1_IN_5 => UNWINDOWED_978 ,
										MUX_10_1_IN_6 => UNWINDOWED_915 ,
										MUX_10_1_IN_7 => UNWINDOWED_915 ,
										MUX_10_1_IN_8 => UNWINDOWED_915 ,
										MUX_10_1_IN_9 => UNWINDOWED_915 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_969
									);
MUX_REORD_UNIT_970 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_970 ,
										MUX_10_1_IN_1 => UNWINDOWED_969 ,
										MUX_10_1_IN_2 => UNWINDOWED_972 ,
										MUX_10_1_IN_3 => UNWINDOWED_965 ,
										MUX_10_1_IN_4 => UNWINDOWED_980 ,
										MUX_10_1_IN_5 => UNWINDOWED_980 ,
										MUX_10_1_IN_6 => UNWINDOWED_917 ,
										MUX_10_1_IN_7 => UNWINDOWED_917 ,
										MUX_10_1_IN_8 => UNWINDOWED_917 ,
										MUX_10_1_IN_9 => UNWINDOWED_917 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_970
									);
MUX_REORD_UNIT_971 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_971 ,
										MUX_10_1_IN_1 => UNWINDOWED_971 ,
										MUX_10_1_IN_2 => UNWINDOWED_974 ,
										MUX_10_1_IN_3 => UNWINDOWED_967 ,
										MUX_10_1_IN_4 => UNWINDOWED_982 ,
										MUX_10_1_IN_5 => UNWINDOWED_982 ,
										MUX_10_1_IN_6 => UNWINDOWED_919 ,
										MUX_10_1_IN_7 => UNWINDOWED_919 ,
										MUX_10_1_IN_8 => UNWINDOWED_919 ,
										MUX_10_1_IN_9 => UNWINDOWED_919 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_971
									);
MUX_REORD_UNIT_972 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_972 ,
										MUX_10_1_IN_1 => UNWINDOWED_972 ,
										MUX_10_1_IN_2 => UNWINDOWED_969 ,
										MUX_10_1_IN_3 => UNWINDOWED_969 ,
										MUX_10_1_IN_4 => UNWINDOWED_984 ,
										MUX_10_1_IN_5 => UNWINDOWED_984 ,
										MUX_10_1_IN_6 => UNWINDOWED_921 ,
										MUX_10_1_IN_7 => UNWINDOWED_921 ,
										MUX_10_1_IN_8 => UNWINDOWED_921 ,
										MUX_10_1_IN_9 => UNWINDOWED_921 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_972
									);
MUX_REORD_UNIT_973 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_973 ,
										MUX_10_1_IN_1 => UNWINDOWED_974 ,
										MUX_10_1_IN_2 => UNWINDOWED_971 ,
										MUX_10_1_IN_3 => UNWINDOWED_971 ,
										MUX_10_1_IN_4 => UNWINDOWED_986 ,
										MUX_10_1_IN_5 => UNWINDOWED_986 ,
										MUX_10_1_IN_6 => UNWINDOWED_923 ,
										MUX_10_1_IN_7 => UNWINDOWED_923 ,
										MUX_10_1_IN_8 => UNWINDOWED_923 ,
										MUX_10_1_IN_9 => UNWINDOWED_923 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_973
									);
MUX_REORD_UNIT_974 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_974 ,
										MUX_10_1_IN_1 => UNWINDOWED_973 ,
										MUX_10_1_IN_2 => UNWINDOWED_973 ,
										MUX_10_1_IN_3 => UNWINDOWED_973 ,
										MUX_10_1_IN_4 => UNWINDOWED_988 ,
										MUX_10_1_IN_5 => UNWINDOWED_988 ,
										MUX_10_1_IN_6 => UNWINDOWED_925 ,
										MUX_10_1_IN_7 => UNWINDOWED_925 ,
										MUX_10_1_IN_8 => UNWINDOWED_925 ,
										MUX_10_1_IN_9 => UNWINDOWED_925 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_974
									);
MUX_REORD_UNIT_975 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_975 ,
										MUX_10_1_IN_1 => UNWINDOWED_975 ,
										MUX_10_1_IN_2 => UNWINDOWED_975 ,
										MUX_10_1_IN_3 => UNWINDOWED_975 ,
										MUX_10_1_IN_4 => UNWINDOWED_990 ,
										MUX_10_1_IN_5 => UNWINDOWED_990 ,
										MUX_10_1_IN_6 => UNWINDOWED_927 ,
										MUX_10_1_IN_7 => UNWINDOWED_927 ,
										MUX_10_1_IN_8 => UNWINDOWED_927 ,
										MUX_10_1_IN_9 => UNWINDOWED_927 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_975
									);
MUX_REORD_UNIT_976 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_976 ,
										MUX_10_1_IN_1 => UNWINDOWED_976 ,
										MUX_10_1_IN_2 => UNWINDOWED_976 ,
										MUX_10_1_IN_3 => UNWINDOWED_976 ,
										MUX_10_1_IN_4 => UNWINDOWED_961 ,
										MUX_10_1_IN_5 => UNWINDOWED_992 ,
										MUX_10_1_IN_6 => UNWINDOWED_929 ,
										MUX_10_1_IN_7 => UNWINDOWED_929 ,
										MUX_10_1_IN_8 => UNWINDOWED_929 ,
										MUX_10_1_IN_9 => UNWINDOWED_929 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_976
									);
MUX_REORD_UNIT_977 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_977 ,
										MUX_10_1_IN_1 => UNWINDOWED_978 ,
										MUX_10_1_IN_2 => UNWINDOWED_978 ,
										MUX_10_1_IN_3 => UNWINDOWED_978 ,
										MUX_10_1_IN_4 => UNWINDOWED_963 ,
										MUX_10_1_IN_5 => UNWINDOWED_994 ,
										MUX_10_1_IN_6 => UNWINDOWED_931 ,
										MUX_10_1_IN_7 => UNWINDOWED_931 ,
										MUX_10_1_IN_8 => UNWINDOWED_931 ,
										MUX_10_1_IN_9 => UNWINDOWED_931 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_977
									);
MUX_REORD_UNIT_978 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_978 ,
										MUX_10_1_IN_1 => UNWINDOWED_977 ,
										MUX_10_1_IN_2 => UNWINDOWED_980 ,
										MUX_10_1_IN_3 => UNWINDOWED_980 ,
										MUX_10_1_IN_4 => UNWINDOWED_965 ,
										MUX_10_1_IN_5 => UNWINDOWED_996 ,
										MUX_10_1_IN_6 => UNWINDOWED_933 ,
										MUX_10_1_IN_7 => UNWINDOWED_933 ,
										MUX_10_1_IN_8 => UNWINDOWED_933 ,
										MUX_10_1_IN_9 => UNWINDOWED_933 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_978
									);
MUX_REORD_UNIT_979 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_979 ,
										MUX_10_1_IN_1 => UNWINDOWED_979 ,
										MUX_10_1_IN_2 => UNWINDOWED_982 ,
										MUX_10_1_IN_3 => UNWINDOWED_982 ,
										MUX_10_1_IN_4 => UNWINDOWED_967 ,
										MUX_10_1_IN_5 => UNWINDOWED_998 ,
										MUX_10_1_IN_6 => UNWINDOWED_935 ,
										MUX_10_1_IN_7 => UNWINDOWED_935 ,
										MUX_10_1_IN_8 => UNWINDOWED_935 ,
										MUX_10_1_IN_9 => UNWINDOWED_935 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_979
									);
MUX_REORD_UNIT_980 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_980 ,
										MUX_10_1_IN_1 => UNWINDOWED_980 ,
										MUX_10_1_IN_2 => UNWINDOWED_977 ,
										MUX_10_1_IN_3 => UNWINDOWED_984 ,
										MUX_10_1_IN_4 => UNWINDOWED_969 ,
										MUX_10_1_IN_5 => UNWINDOWED_1000 ,
										MUX_10_1_IN_6 => UNWINDOWED_937 ,
										MUX_10_1_IN_7 => UNWINDOWED_937 ,
										MUX_10_1_IN_8 => UNWINDOWED_937 ,
										MUX_10_1_IN_9 => UNWINDOWED_937 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_980
									);
MUX_REORD_UNIT_981 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_981 ,
										MUX_10_1_IN_1 => UNWINDOWED_982 ,
										MUX_10_1_IN_2 => UNWINDOWED_979 ,
										MUX_10_1_IN_3 => UNWINDOWED_986 ,
										MUX_10_1_IN_4 => UNWINDOWED_971 ,
										MUX_10_1_IN_5 => UNWINDOWED_1002 ,
										MUX_10_1_IN_6 => UNWINDOWED_939 ,
										MUX_10_1_IN_7 => UNWINDOWED_939 ,
										MUX_10_1_IN_8 => UNWINDOWED_939 ,
										MUX_10_1_IN_9 => UNWINDOWED_939 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_981
									);
MUX_REORD_UNIT_982 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_982 ,
										MUX_10_1_IN_1 => UNWINDOWED_981 ,
										MUX_10_1_IN_2 => UNWINDOWED_981 ,
										MUX_10_1_IN_3 => UNWINDOWED_988 ,
										MUX_10_1_IN_4 => UNWINDOWED_973 ,
										MUX_10_1_IN_5 => UNWINDOWED_1004 ,
										MUX_10_1_IN_6 => UNWINDOWED_941 ,
										MUX_10_1_IN_7 => UNWINDOWED_941 ,
										MUX_10_1_IN_8 => UNWINDOWED_941 ,
										MUX_10_1_IN_9 => UNWINDOWED_941 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_982
									);
MUX_REORD_UNIT_983 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_983 ,
										MUX_10_1_IN_1 => UNWINDOWED_983 ,
										MUX_10_1_IN_2 => UNWINDOWED_983 ,
										MUX_10_1_IN_3 => UNWINDOWED_990 ,
										MUX_10_1_IN_4 => UNWINDOWED_975 ,
										MUX_10_1_IN_5 => UNWINDOWED_1006 ,
										MUX_10_1_IN_6 => UNWINDOWED_943 ,
										MUX_10_1_IN_7 => UNWINDOWED_943 ,
										MUX_10_1_IN_8 => UNWINDOWED_943 ,
										MUX_10_1_IN_9 => UNWINDOWED_943 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_983
									);
MUX_REORD_UNIT_984 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_984 ,
										MUX_10_1_IN_1 => UNWINDOWED_984 ,
										MUX_10_1_IN_2 => UNWINDOWED_984 ,
										MUX_10_1_IN_3 => UNWINDOWED_977 ,
										MUX_10_1_IN_4 => UNWINDOWED_977 ,
										MUX_10_1_IN_5 => UNWINDOWED_1008 ,
										MUX_10_1_IN_6 => UNWINDOWED_945 ,
										MUX_10_1_IN_7 => UNWINDOWED_945 ,
										MUX_10_1_IN_8 => UNWINDOWED_945 ,
										MUX_10_1_IN_9 => UNWINDOWED_945 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_984
									);
MUX_REORD_UNIT_985 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_985 ,
										MUX_10_1_IN_1 => UNWINDOWED_986 ,
										MUX_10_1_IN_2 => UNWINDOWED_986 ,
										MUX_10_1_IN_3 => UNWINDOWED_979 ,
										MUX_10_1_IN_4 => UNWINDOWED_979 ,
										MUX_10_1_IN_5 => UNWINDOWED_1010 ,
										MUX_10_1_IN_6 => UNWINDOWED_947 ,
										MUX_10_1_IN_7 => UNWINDOWED_947 ,
										MUX_10_1_IN_8 => UNWINDOWED_947 ,
										MUX_10_1_IN_9 => UNWINDOWED_947 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_985
									);
MUX_REORD_UNIT_986 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_986 ,
										MUX_10_1_IN_1 => UNWINDOWED_985 ,
										MUX_10_1_IN_2 => UNWINDOWED_988 ,
										MUX_10_1_IN_3 => UNWINDOWED_981 ,
										MUX_10_1_IN_4 => UNWINDOWED_981 ,
										MUX_10_1_IN_5 => UNWINDOWED_1012 ,
										MUX_10_1_IN_6 => UNWINDOWED_949 ,
										MUX_10_1_IN_7 => UNWINDOWED_949 ,
										MUX_10_1_IN_8 => UNWINDOWED_949 ,
										MUX_10_1_IN_9 => UNWINDOWED_949 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_986
									);
MUX_REORD_UNIT_987 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_987 ,
										MUX_10_1_IN_1 => UNWINDOWED_987 ,
										MUX_10_1_IN_2 => UNWINDOWED_990 ,
										MUX_10_1_IN_3 => UNWINDOWED_983 ,
										MUX_10_1_IN_4 => UNWINDOWED_983 ,
										MUX_10_1_IN_5 => UNWINDOWED_1014 ,
										MUX_10_1_IN_6 => UNWINDOWED_951 ,
										MUX_10_1_IN_7 => UNWINDOWED_951 ,
										MUX_10_1_IN_8 => UNWINDOWED_951 ,
										MUX_10_1_IN_9 => UNWINDOWED_951 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_987
									);
MUX_REORD_UNIT_988 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_988 ,
										MUX_10_1_IN_1 => UNWINDOWED_988 ,
										MUX_10_1_IN_2 => UNWINDOWED_985 ,
										MUX_10_1_IN_3 => UNWINDOWED_985 ,
										MUX_10_1_IN_4 => UNWINDOWED_985 ,
										MUX_10_1_IN_5 => UNWINDOWED_1016 ,
										MUX_10_1_IN_6 => UNWINDOWED_953 ,
										MUX_10_1_IN_7 => UNWINDOWED_953 ,
										MUX_10_1_IN_8 => UNWINDOWED_953 ,
										MUX_10_1_IN_9 => UNWINDOWED_953 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_988
									);
MUX_REORD_UNIT_989 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_989 ,
										MUX_10_1_IN_1 => UNWINDOWED_990 ,
										MUX_10_1_IN_2 => UNWINDOWED_987 ,
										MUX_10_1_IN_3 => UNWINDOWED_987 ,
										MUX_10_1_IN_4 => UNWINDOWED_987 ,
										MUX_10_1_IN_5 => UNWINDOWED_1018 ,
										MUX_10_1_IN_6 => UNWINDOWED_955 ,
										MUX_10_1_IN_7 => UNWINDOWED_955 ,
										MUX_10_1_IN_8 => UNWINDOWED_955 ,
										MUX_10_1_IN_9 => UNWINDOWED_955 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_989
									);
MUX_REORD_UNIT_990 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_990 ,
										MUX_10_1_IN_1 => UNWINDOWED_989 ,
										MUX_10_1_IN_2 => UNWINDOWED_989 ,
										MUX_10_1_IN_3 => UNWINDOWED_989 ,
										MUX_10_1_IN_4 => UNWINDOWED_989 ,
										MUX_10_1_IN_5 => UNWINDOWED_1020 ,
										MUX_10_1_IN_6 => UNWINDOWED_957 ,
										MUX_10_1_IN_7 => UNWINDOWED_957 ,
										MUX_10_1_IN_8 => UNWINDOWED_957 ,
										MUX_10_1_IN_9 => UNWINDOWED_957 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_990
									);
MUX_REORD_UNIT_991 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_991 ,
										MUX_10_1_IN_1 => UNWINDOWED_991 ,
										MUX_10_1_IN_2 => UNWINDOWED_991 ,
										MUX_10_1_IN_3 => UNWINDOWED_991 ,
										MUX_10_1_IN_4 => UNWINDOWED_991 ,
										MUX_10_1_IN_5 => UNWINDOWED_1022 ,
										MUX_10_1_IN_6 => UNWINDOWED_959 ,
										MUX_10_1_IN_7 => UNWINDOWED_959 ,
										MUX_10_1_IN_8 => UNWINDOWED_959 ,
										MUX_10_1_IN_9 => UNWINDOWED_959 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_991
									);
MUX_REORD_UNIT_992 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_992 ,
										MUX_10_1_IN_1 => UNWINDOWED_992 ,
										MUX_10_1_IN_2 => UNWINDOWED_992 ,
										MUX_10_1_IN_3 => UNWINDOWED_992 ,
										MUX_10_1_IN_4 => UNWINDOWED_992 ,
										MUX_10_1_IN_5 => UNWINDOWED_961 ,
										MUX_10_1_IN_6 => UNWINDOWED_961 ,
										MUX_10_1_IN_7 => UNWINDOWED_961 ,
										MUX_10_1_IN_8 => UNWINDOWED_961 ,
										MUX_10_1_IN_9 => UNWINDOWED_961 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_992
									);
MUX_REORD_UNIT_993 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_993 ,
										MUX_10_1_IN_1 => UNWINDOWED_994 ,
										MUX_10_1_IN_2 => UNWINDOWED_994 ,
										MUX_10_1_IN_3 => UNWINDOWED_994 ,
										MUX_10_1_IN_4 => UNWINDOWED_994 ,
										MUX_10_1_IN_5 => UNWINDOWED_963 ,
										MUX_10_1_IN_6 => UNWINDOWED_963 ,
										MUX_10_1_IN_7 => UNWINDOWED_963 ,
										MUX_10_1_IN_8 => UNWINDOWED_963 ,
										MUX_10_1_IN_9 => UNWINDOWED_963 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_993
									);
MUX_REORD_UNIT_994 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_994 ,
										MUX_10_1_IN_1 => UNWINDOWED_993 ,
										MUX_10_1_IN_2 => UNWINDOWED_996 ,
										MUX_10_1_IN_3 => UNWINDOWED_996 ,
										MUX_10_1_IN_4 => UNWINDOWED_996 ,
										MUX_10_1_IN_5 => UNWINDOWED_965 ,
										MUX_10_1_IN_6 => UNWINDOWED_965 ,
										MUX_10_1_IN_7 => UNWINDOWED_965 ,
										MUX_10_1_IN_8 => UNWINDOWED_965 ,
										MUX_10_1_IN_9 => UNWINDOWED_965 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_994
									);
MUX_REORD_UNIT_995 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_995 ,
										MUX_10_1_IN_1 => UNWINDOWED_995 ,
										MUX_10_1_IN_2 => UNWINDOWED_998 ,
										MUX_10_1_IN_3 => UNWINDOWED_998 ,
										MUX_10_1_IN_4 => UNWINDOWED_998 ,
										MUX_10_1_IN_5 => UNWINDOWED_967 ,
										MUX_10_1_IN_6 => UNWINDOWED_967 ,
										MUX_10_1_IN_7 => UNWINDOWED_967 ,
										MUX_10_1_IN_8 => UNWINDOWED_967 ,
										MUX_10_1_IN_9 => UNWINDOWED_967 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_995
									);
MUX_REORD_UNIT_996 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_996 ,
										MUX_10_1_IN_1 => UNWINDOWED_996 ,
										MUX_10_1_IN_2 => UNWINDOWED_993 ,
										MUX_10_1_IN_3 => UNWINDOWED_1000 ,
										MUX_10_1_IN_4 => UNWINDOWED_1000 ,
										MUX_10_1_IN_5 => UNWINDOWED_969 ,
										MUX_10_1_IN_6 => UNWINDOWED_969 ,
										MUX_10_1_IN_7 => UNWINDOWED_969 ,
										MUX_10_1_IN_8 => UNWINDOWED_969 ,
										MUX_10_1_IN_9 => UNWINDOWED_969 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_996
									);
MUX_REORD_UNIT_997 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_997 ,
										MUX_10_1_IN_1 => UNWINDOWED_998 ,
										MUX_10_1_IN_2 => UNWINDOWED_995 ,
										MUX_10_1_IN_3 => UNWINDOWED_1002 ,
										MUX_10_1_IN_4 => UNWINDOWED_1002 ,
										MUX_10_1_IN_5 => UNWINDOWED_971 ,
										MUX_10_1_IN_6 => UNWINDOWED_971 ,
										MUX_10_1_IN_7 => UNWINDOWED_971 ,
										MUX_10_1_IN_8 => UNWINDOWED_971 ,
										MUX_10_1_IN_9 => UNWINDOWED_971 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_997
									);
MUX_REORD_UNIT_998 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_998 ,
										MUX_10_1_IN_1 => UNWINDOWED_997 ,
										MUX_10_1_IN_2 => UNWINDOWED_997 ,
										MUX_10_1_IN_3 => UNWINDOWED_1004 ,
										MUX_10_1_IN_4 => UNWINDOWED_1004 ,
										MUX_10_1_IN_5 => UNWINDOWED_973 ,
										MUX_10_1_IN_6 => UNWINDOWED_973 ,
										MUX_10_1_IN_7 => UNWINDOWED_973 ,
										MUX_10_1_IN_8 => UNWINDOWED_973 ,
										MUX_10_1_IN_9 => UNWINDOWED_973 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_998
									);
MUX_REORD_UNIT_999 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_999 ,
										MUX_10_1_IN_1 => UNWINDOWED_999 ,
										MUX_10_1_IN_2 => UNWINDOWED_999 ,
										MUX_10_1_IN_3 => UNWINDOWED_1006 ,
										MUX_10_1_IN_4 => UNWINDOWED_1006 ,
										MUX_10_1_IN_5 => UNWINDOWED_975 ,
										MUX_10_1_IN_6 => UNWINDOWED_975 ,
										MUX_10_1_IN_7 => UNWINDOWED_975 ,
										MUX_10_1_IN_8 => UNWINDOWED_975 ,
										MUX_10_1_IN_9 => UNWINDOWED_975 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_999
									);
MUX_REORD_UNIT_1000 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1000 ,
										MUX_10_1_IN_1 => UNWINDOWED_1000 ,
										MUX_10_1_IN_2 => UNWINDOWED_1000 ,
										MUX_10_1_IN_3 => UNWINDOWED_993 ,
										MUX_10_1_IN_4 => UNWINDOWED_1008 ,
										MUX_10_1_IN_5 => UNWINDOWED_977 ,
										MUX_10_1_IN_6 => UNWINDOWED_977 ,
										MUX_10_1_IN_7 => UNWINDOWED_977 ,
										MUX_10_1_IN_8 => UNWINDOWED_977 ,
										MUX_10_1_IN_9 => UNWINDOWED_977 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1000
									);
MUX_REORD_UNIT_1001 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1001 ,
										MUX_10_1_IN_1 => UNWINDOWED_1002 ,
										MUX_10_1_IN_2 => UNWINDOWED_1002 ,
										MUX_10_1_IN_3 => UNWINDOWED_995 ,
										MUX_10_1_IN_4 => UNWINDOWED_1010 ,
										MUX_10_1_IN_5 => UNWINDOWED_979 ,
										MUX_10_1_IN_6 => UNWINDOWED_979 ,
										MUX_10_1_IN_7 => UNWINDOWED_979 ,
										MUX_10_1_IN_8 => UNWINDOWED_979 ,
										MUX_10_1_IN_9 => UNWINDOWED_979 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1001
									);
MUX_REORD_UNIT_1002 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1002 ,
										MUX_10_1_IN_1 => UNWINDOWED_1001 ,
										MUX_10_1_IN_2 => UNWINDOWED_1004 ,
										MUX_10_1_IN_3 => UNWINDOWED_997 ,
										MUX_10_1_IN_4 => UNWINDOWED_1012 ,
										MUX_10_1_IN_5 => UNWINDOWED_981 ,
										MUX_10_1_IN_6 => UNWINDOWED_981 ,
										MUX_10_1_IN_7 => UNWINDOWED_981 ,
										MUX_10_1_IN_8 => UNWINDOWED_981 ,
										MUX_10_1_IN_9 => UNWINDOWED_981 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1002
									);
MUX_REORD_UNIT_1003 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1003 ,
										MUX_10_1_IN_1 => UNWINDOWED_1003 ,
										MUX_10_1_IN_2 => UNWINDOWED_1006 ,
										MUX_10_1_IN_3 => UNWINDOWED_999 ,
										MUX_10_1_IN_4 => UNWINDOWED_1014 ,
										MUX_10_1_IN_5 => UNWINDOWED_983 ,
										MUX_10_1_IN_6 => UNWINDOWED_983 ,
										MUX_10_1_IN_7 => UNWINDOWED_983 ,
										MUX_10_1_IN_8 => UNWINDOWED_983 ,
										MUX_10_1_IN_9 => UNWINDOWED_983 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1003
									);
MUX_REORD_UNIT_1004 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1004 ,
										MUX_10_1_IN_1 => UNWINDOWED_1004 ,
										MUX_10_1_IN_2 => UNWINDOWED_1001 ,
										MUX_10_1_IN_3 => UNWINDOWED_1001 ,
										MUX_10_1_IN_4 => UNWINDOWED_1016 ,
										MUX_10_1_IN_5 => UNWINDOWED_985 ,
										MUX_10_1_IN_6 => UNWINDOWED_985 ,
										MUX_10_1_IN_7 => UNWINDOWED_985 ,
										MUX_10_1_IN_8 => UNWINDOWED_985 ,
										MUX_10_1_IN_9 => UNWINDOWED_985 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1004
									);
MUX_REORD_UNIT_1005 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1005 ,
										MUX_10_1_IN_1 => UNWINDOWED_1006 ,
										MUX_10_1_IN_2 => UNWINDOWED_1003 ,
										MUX_10_1_IN_3 => UNWINDOWED_1003 ,
										MUX_10_1_IN_4 => UNWINDOWED_1018 ,
										MUX_10_1_IN_5 => UNWINDOWED_987 ,
										MUX_10_1_IN_6 => UNWINDOWED_987 ,
										MUX_10_1_IN_7 => UNWINDOWED_987 ,
										MUX_10_1_IN_8 => UNWINDOWED_987 ,
										MUX_10_1_IN_9 => UNWINDOWED_987 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1005
									);
MUX_REORD_UNIT_1006 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1006 ,
										MUX_10_1_IN_1 => UNWINDOWED_1005 ,
										MUX_10_1_IN_2 => UNWINDOWED_1005 ,
										MUX_10_1_IN_3 => UNWINDOWED_1005 ,
										MUX_10_1_IN_4 => UNWINDOWED_1020 ,
										MUX_10_1_IN_5 => UNWINDOWED_989 ,
										MUX_10_1_IN_6 => UNWINDOWED_989 ,
										MUX_10_1_IN_7 => UNWINDOWED_989 ,
										MUX_10_1_IN_8 => UNWINDOWED_989 ,
										MUX_10_1_IN_9 => UNWINDOWED_989 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1006
									);
MUX_REORD_UNIT_1007 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1007 ,
										MUX_10_1_IN_1 => UNWINDOWED_1007 ,
										MUX_10_1_IN_2 => UNWINDOWED_1007 ,
										MUX_10_1_IN_3 => UNWINDOWED_1007 ,
										MUX_10_1_IN_4 => UNWINDOWED_1022 ,
										MUX_10_1_IN_5 => UNWINDOWED_991 ,
										MUX_10_1_IN_6 => UNWINDOWED_991 ,
										MUX_10_1_IN_7 => UNWINDOWED_991 ,
										MUX_10_1_IN_8 => UNWINDOWED_991 ,
										MUX_10_1_IN_9 => UNWINDOWED_991 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1007
									);
MUX_REORD_UNIT_1008 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1008 ,
										MUX_10_1_IN_1 => UNWINDOWED_1008 ,
										MUX_10_1_IN_2 => UNWINDOWED_1008 ,
										MUX_10_1_IN_3 => UNWINDOWED_1008 ,
										MUX_10_1_IN_4 => UNWINDOWED_993 ,
										MUX_10_1_IN_5 => UNWINDOWED_993 ,
										MUX_10_1_IN_6 => UNWINDOWED_993 ,
										MUX_10_1_IN_7 => UNWINDOWED_993 ,
										MUX_10_1_IN_8 => UNWINDOWED_993 ,
										MUX_10_1_IN_9 => UNWINDOWED_993 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1008
									);
MUX_REORD_UNIT_1009 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1009 ,
										MUX_10_1_IN_1 => UNWINDOWED_1010 ,
										MUX_10_1_IN_2 => UNWINDOWED_1010 ,
										MUX_10_1_IN_3 => UNWINDOWED_1010 ,
										MUX_10_1_IN_4 => UNWINDOWED_995 ,
										MUX_10_1_IN_5 => UNWINDOWED_995 ,
										MUX_10_1_IN_6 => UNWINDOWED_995 ,
										MUX_10_1_IN_7 => UNWINDOWED_995 ,
										MUX_10_1_IN_8 => UNWINDOWED_995 ,
										MUX_10_1_IN_9 => UNWINDOWED_995 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1009
									);
MUX_REORD_UNIT_1010 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1010 ,
										MUX_10_1_IN_1 => UNWINDOWED_1009 ,
										MUX_10_1_IN_2 => UNWINDOWED_1012 ,
										MUX_10_1_IN_3 => UNWINDOWED_1012 ,
										MUX_10_1_IN_4 => UNWINDOWED_997 ,
										MUX_10_1_IN_5 => UNWINDOWED_997 ,
										MUX_10_1_IN_6 => UNWINDOWED_997 ,
										MUX_10_1_IN_7 => UNWINDOWED_997 ,
										MUX_10_1_IN_8 => UNWINDOWED_997 ,
										MUX_10_1_IN_9 => UNWINDOWED_997 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1010
									);
MUX_REORD_UNIT_1011 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1011 ,
										MUX_10_1_IN_1 => UNWINDOWED_1011 ,
										MUX_10_1_IN_2 => UNWINDOWED_1014 ,
										MUX_10_1_IN_3 => UNWINDOWED_1014 ,
										MUX_10_1_IN_4 => UNWINDOWED_999 ,
										MUX_10_1_IN_5 => UNWINDOWED_999 ,
										MUX_10_1_IN_6 => UNWINDOWED_999 ,
										MUX_10_1_IN_7 => UNWINDOWED_999 ,
										MUX_10_1_IN_8 => UNWINDOWED_999 ,
										MUX_10_1_IN_9 => UNWINDOWED_999 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1011
									);
MUX_REORD_UNIT_1012 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1012 ,
										MUX_10_1_IN_1 => UNWINDOWED_1012 ,
										MUX_10_1_IN_2 => UNWINDOWED_1009 ,
										MUX_10_1_IN_3 => UNWINDOWED_1016 ,
										MUX_10_1_IN_4 => UNWINDOWED_1001 ,
										MUX_10_1_IN_5 => UNWINDOWED_1001 ,
										MUX_10_1_IN_6 => UNWINDOWED_1001 ,
										MUX_10_1_IN_7 => UNWINDOWED_1001 ,
										MUX_10_1_IN_8 => UNWINDOWED_1001 ,
										MUX_10_1_IN_9 => UNWINDOWED_1001 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1012
									);
MUX_REORD_UNIT_1013 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1013 ,
										MUX_10_1_IN_1 => UNWINDOWED_1014 ,
										MUX_10_1_IN_2 => UNWINDOWED_1011 ,
										MUX_10_1_IN_3 => UNWINDOWED_1018 ,
										MUX_10_1_IN_4 => UNWINDOWED_1003 ,
										MUX_10_1_IN_5 => UNWINDOWED_1003 ,
										MUX_10_1_IN_6 => UNWINDOWED_1003 ,
										MUX_10_1_IN_7 => UNWINDOWED_1003 ,
										MUX_10_1_IN_8 => UNWINDOWED_1003 ,
										MUX_10_1_IN_9 => UNWINDOWED_1003 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1013
									);
MUX_REORD_UNIT_1014 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1014 ,
										MUX_10_1_IN_1 => UNWINDOWED_1013 ,
										MUX_10_1_IN_2 => UNWINDOWED_1013 ,
										MUX_10_1_IN_3 => UNWINDOWED_1020 ,
										MUX_10_1_IN_4 => UNWINDOWED_1005 ,
										MUX_10_1_IN_5 => UNWINDOWED_1005 ,
										MUX_10_1_IN_6 => UNWINDOWED_1005 ,
										MUX_10_1_IN_7 => UNWINDOWED_1005 ,
										MUX_10_1_IN_8 => UNWINDOWED_1005 ,
										MUX_10_1_IN_9 => UNWINDOWED_1005 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1014
									);
MUX_REORD_UNIT_1015 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1015 ,
										MUX_10_1_IN_1 => UNWINDOWED_1015 ,
										MUX_10_1_IN_2 => UNWINDOWED_1015 ,
										MUX_10_1_IN_3 => UNWINDOWED_1022 ,
										MUX_10_1_IN_4 => UNWINDOWED_1007 ,
										MUX_10_1_IN_5 => UNWINDOWED_1007 ,
										MUX_10_1_IN_6 => UNWINDOWED_1007 ,
										MUX_10_1_IN_7 => UNWINDOWED_1007 ,
										MUX_10_1_IN_8 => UNWINDOWED_1007 ,
										MUX_10_1_IN_9 => UNWINDOWED_1007 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1015
									);
MUX_REORD_UNIT_1016 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1016 ,
										MUX_10_1_IN_1 => UNWINDOWED_1016 ,
										MUX_10_1_IN_2 => UNWINDOWED_1016 ,
										MUX_10_1_IN_3 => UNWINDOWED_1009 ,
										MUX_10_1_IN_4 => UNWINDOWED_1009 ,
										MUX_10_1_IN_5 => UNWINDOWED_1009 ,
										MUX_10_1_IN_6 => UNWINDOWED_1009 ,
										MUX_10_1_IN_7 => UNWINDOWED_1009 ,
										MUX_10_1_IN_8 => UNWINDOWED_1009 ,
										MUX_10_1_IN_9 => UNWINDOWED_1009 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1016
									);
MUX_REORD_UNIT_1017 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1017 ,
										MUX_10_1_IN_1 => UNWINDOWED_1018 ,
										MUX_10_1_IN_2 => UNWINDOWED_1018 ,
										MUX_10_1_IN_3 => UNWINDOWED_1011 ,
										MUX_10_1_IN_4 => UNWINDOWED_1011 ,
										MUX_10_1_IN_5 => UNWINDOWED_1011 ,
										MUX_10_1_IN_6 => UNWINDOWED_1011 ,
										MUX_10_1_IN_7 => UNWINDOWED_1011 ,
										MUX_10_1_IN_8 => UNWINDOWED_1011 ,
										MUX_10_1_IN_9 => UNWINDOWED_1011 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1017
									);
MUX_REORD_UNIT_1018 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1018 ,
										MUX_10_1_IN_1 => UNWINDOWED_1017 ,
										MUX_10_1_IN_2 => UNWINDOWED_1020 ,
										MUX_10_1_IN_3 => UNWINDOWED_1013 ,
										MUX_10_1_IN_4 => UNWINDOWED_1013 ,
										MUX_10_1_IN_5 => UNWINDOWED_1013 ,
										MUX_10_1_IN_6 => UNWINDOWED_1013 ,
										MUX_10_1_IN_7 => UNWINDOWED_1013 ,
										MUX_10_1_IN_8 => UNWINDOWED_1013 ,
										MUX_10_1_IN_9 => UNWINDOWED_1013 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1018
									);
MUX_REORD_UNIT_1019 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1019 ,
										MUX_10_1_IN_1 => UNWINDOWED_1019 ,
										MUX_10_1_IN_2 => UNWINDOWED_1022 ,
										MUX_10_1_IN_3 => UNWINDOWED_1015 ,
										MUX_10_1_IN_4 => UNWINDOWED_1015 ,
										MUX_10_1_IN_5 => UNWINDOWED_1015 ,
										MUX_10_1_IN_6 => UNWINDOWED_1015 ,
										MUX_10_1_IN_7 => UNWINDOWED_1015 ,
										MUX_10_1_IN_8 => UNWINDOWED_1015 ,
										MUX_10_1_IN_9 => UNWINDOWED_1015 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1019
									);
MUX_REORD_UNIT_1020 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1020 ,
										MUX_10_1_IN_1 => UNWINDOWED_1020 ,
										MUX_10_1_IN_2 => UNWINDOWED_1017 ,
										MUX_10_1_IN_3 => UNWINDOWED_1017 ,
										MUX_10_1_IN_4 => UNWINDOWED_1017 ,
										MUX_10_1_IN_5 => UNWINDOWED_1017 ,
										MUX_10_1_IN_6 => UNWINDOWED_1017 ,
										MUX_10_1_IN_7 => UNWINDOWED_1017 ,
										MUX_10_1_IN_8 => UNWINDOWED_1017 ,
										MUX_10_1_IN_9 => UNWINDOWED_1017 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1020
									);
MUX_REORD_UNIT_1021 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1021 ,
										MUX_10_1_IN_1 => UNWINDOWED_1022 ,
										MUX_10_1_IN_2 => UNWINDOWED_1019 ,
										MUX_10_1_IN_3 => UNWINDOWED_1019 ,
										MUX_10_1_IN_4 => UNWINDOWED_1019 ,
										MUX_10_1_IN_5 => UNWINDOWED_1019 ,
										MUX_10_1_IN_6 => UNWINDOWED_1019 ,
										MUX_10_1_IN_7 => UNWINDOWED_1019 ,
										MUX_10_1_IN_8 => UNWINDOWED_1019 ,
										MUX_10_1_IN_9 => UNWINDOWED_1019 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1021
									);
MUX_REORD_UNIT_1022 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1022 ,
										MUX_10_1_IN_1 => UNWINDOWED_1021 ,
										MUX_10_1_IN_2 => UNWINDOWED_1021 ,
										MUX_10_1_IN_3 => UNWINDOWED_1021 ,
										MUX_10_1_IN_4 => UNWINDOWED_1021 ,
										MUX_10_1_IN_5 => UNWINDOWED_1021 ,
										MUX_10_1_IN_6 => UNWINDOWED_1021 ,
										MUX_10_1_IN_7 => UNWINDOWED_1021 ,
										MUX_10_1_IN_8 => UNWINDOWED_1021 ,
										MUX_10_1_IN_9 => UNWINDOWED_1021 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1022
									);
MUX_REORD_UNIT_1023 : multiplexer_10_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_10_1_IN_0 => UNWINDOWED_1023 ,
										MUX_10_1_IN_1 => UNWINDOWED_1023 ,
										MUX_10_1_IN_2 => UNWINDOWED_1023 ,
										MUX_10_1_IN_3 => UNWINDOWED_1023 ,
										MUX_10_1_IN_4 => UNWINDOWED_1023 ,
										MUX_10_1_IN_5 => UNWINDOWED_1023 ,
										MUX_10_1_IN_6 => UNWINDOWED_1023 ,
										MUX_10_1_IN_7 => UNWINDOWED_1023 ,
										MUX_10_1_IN_8 => UNWINDOWED_1023 ,
										MUX_10_1_IN_9 => UNWINDOWED_1023 ,
				                    			MUX_10_1_IN_SEL => QEP_N_10_W_0_S_0_IN_QTGT ,
										MUX_10_1_OUT_RES => TO_STATE_REG_1023
									);

MUX_OUTPUT_SELECTION : multiplexer_1024_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_1024_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_1024_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_1024_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_1024_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_1024_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_1024_1_IN_5 => FROM_STATE_REG_5 ,
										MUX_1024_1_IN_6 => FROM_STATE_REG_6 ,
										MUX_1024_1_IN_7 => FROM_STATE_REG_7 ,
										MUX_1024_1_IN_8 => FROM_STATE_REG_8 ,
										MUX_1024_1_IN_9 => FROM_STATE_REG_9 ,
										MUX_1024_1_IN_10 => FROM_STATE_REG_10 ,
										MUX_1024_1_IN_11 => FROM_STATE_REG_11 ,
										MUX_1024_1_IN_12 => FROM_STATE_REG_12 ,
										MUX_1024_1_IN_13 => FROM_STATE_REG_13 ,
										MUX_1024_1_IN_14 => FROM_STATE_REG_14 ,
										MUX_1024_1_IN_15 => FROM_STATE_REG_15 ,
										MUX_1024_1_IN_16 => FROM_STATE_REG_16 ,
										MUX_1024_1_IN_17 => FROM_STATE_REG_17 ,
										MUX_1024_1_IN_18 => FROM_STATE_REG_18 ,
										MUX_1024_1_IN_19 => FROM_STATE_REG_19 ,
										MUX_1024_1_IN_20 => FROM_STATE_REG_20 ,
										MUX_1024_1_IN_21 => FROM_STATE_REG_21 ,
										MUX_1024_1_IN_22 => FROM_STATE_REG_22 ,
										MUX_1024_1_IN_23 => FROM_STATE_REG_23 ,
										MUX_1024_1_IN_24 => FROM_STATE_REG_24 ,
										MUX_1024_1_IN_25 => FROM_STATE_REG_25 ,
										MUX_1024_1_IN_26 => FROM_STATE_REG_26 ,
										MUX_1024_1_IN_27 => FROM_STATE_REG_27 ,
										MUX_1024_1_IN_28 => FROM_STATE_REG_28 ,
										MUX_1024_1_IN_29 => FROM_STATE_REG_29 ,
										MUX_1024_1_IN_30 => FROM_STATE_REG_30 ,
										MUX_1024_1_IN_31 => FROM_STATE_REG_31 ,
										MUX_1024_1_IN_32 => FROM_STATE_REG_32 ,
										MUX_1024_1_IN_33 => FROM_STATE_REG_33 ,
										MUX_1024_1_IN_34 => FROM_STATE_REG_34 ,
										MUX_1024_1_IN_35 => FROM_STATE_REG_35 ,
										MUX_1024_1_IN_36 => FROM_STATE_REG_36 ,
										MUX_1024_1_IN_37 => FROM_STATE_REG_37 ,
										MUX_1024_1_IN_38 => FROM_STATE_REG_38 ,
										MUX_1024_1_IN_39 => FROM_STATE_REG_39 ,
										MUX_1024_1_IN_40 => FROM_STATE_REG_40 ,
										MUX_1024_1_IN_41 => FROM_STATE_REG_41 ,
										MUX_1024_1_IN_42 => FROM_STATE_REG_42 ,
										MUX_1024_1_IN_43 => FROM_STATE_REG_43 ,
										MUX_1024_1_IN_44 => FROM_STATE_REG_44 ,
										MUX_1024_1_IN_45 => FROM_STATE_REG_45 ,
										MUX_1024_1_IN_46 => FROM_STATE_REG_46 ,
										MUX_1024_1_IN_47 => FROM_STATE_REG_47 ,
										MUX_1024_1_IN_48 => FROM_STATE_REG_48 ,
										MUX_1024_1_IN_49 => FROM_STATE_REG_49 ,
										MUX_1024_1_IN_50 => FROM_STATE_REG_50 ,
										MUX_1024_1_IN_51 => FROM_STATE_REG_51 ,
										MUX_1024_1_IN_52 => FROM_STATE_REG_52 ,
										MUX_1024_1_IN_53 => FROM_STATE_REG_53 ,
										MUX_1024_1_IN_54 => FROM_STATE_REG_54 ,
										MUX_1024_1_IN_55 => FROM_STATE_REG_55 ,
										MUX_1024_1_IN_56 => FROM_STATE_REG_56 ,
										MUX_1024_1_IN_57 => FROM_STATE_REG_57 ,
										MUX_1024_1_IN_58 => FROM_STATE_REG_58 ,
										MUX_1024_1_IN_59 => FROM_STATE_REG_59 ,
										MUX_1024_1_IN_60 => FROM_STATE_REG_60 ,
										MUX_1024_1_IN_61 => FROM_STATE_REG_61 ,
										MUX_1024_1_IN_62 => FROM_STATE_REG_62 ,
										MUX_1024_1_IN_63 => FROM_STATE_REG_63 ,
										MUX_1024_1_IN_64 => FROM_STATE_REG_64 ,
										MUX_1024_1_IN_65 => FROM_STATE_REG_65 ,
										MUX_1024_1_IN_66 => FROM_STATE_REG_66 ,
										MUX_1024_1_IN_67 => FROM_STATE_REG_67 ,
										MUX_1024_1_IN_68 => FROM_STATE_REG_68 ,
										MUX_1024_1_IN_69 => FROM_STATE_REG_69 ,
										MUX_1024_1_IN_70 => FROM_STATE_REG_70 ,
										MUX_1024_1_IN_71 => FROM_STATE_REG_71 ,
										MUX_1024_1_IN_72 => FROM_STATE_REG_72 ,
										MUX_1024_1_IN_73 => FROM_STATE_REG_73 ,
										MUX_1024_1_IN_74 => FROM_STATE_REG_74 ,
										MUX_1024_1_IN_75 => FROM_STATE_REG_75 ,
										MUX_1024_1_IN_76 => FROM_STATE_REG_76 ,
										MUX_1024_1_IN_77 => FROM_STATE_REG_77 ,
										MUX_1024_1_IN_78 => FROM_STATE_REG_78 ,
										MUX_1024_1_IN_79 => FROM_STATE_REG_79 ,
										MUX_1024_1_IN_80 => FROM_STATE_REG_80 ,
										MUX_1024_1_IN_81 => FROM_STATE_REG_81 ,
										MUX_1024_1_IN_82 => FROM_STATE_REG_82 ,
										MUX_1024_1_IN_83 => FROM_STATE_REG_83 ,
										MUX_1024_1_IN_84 => FROM_STATE_REG_84 ,
										MUX_1024_1_IN_85 => FROM_STATE_REG_85 ,
										MUX_1024_1_IN_86 => FROM_STATE_REG_86 ,
										MUX_1024_1_IN_87 => FROM_STATE_REG_87 ,
										MUX_1024_1_IN_88 => FROM_STATE_REG_88 ,
										MUX_1024_1_IN_89 => FROM_STATE_REG_89 ,
										MUX_1024_1_IN_90 => FROM_STATE_REG_90 ,
										MUX_1024_1_IN_91 => FROM_STATE_REG_91 ,
										MUX_1024_1_IN_92 => FROM_STATE_REG_92 ,
										MUX_1024_1_IN_93 => FROM_STATE_REG_93 ,
										MUX_1024_1_IN_94 => FROM_STATE_REG_94 ,
										MUX_1024_1_IN_95 => FROM_STATE_REG_95 ,
										MUX_1024_1_IN_96 => FROM_STATE_REG_96 ,
										MUX_1024_1_IN_97 => FROM_STATE_REG_97 ,
										MUX_1024_1_IN_98 => FROM_STATE_REG_98 ,
										MUX_1024_1_IN_99 => FROM_STATE_REG_99 ,
										MUX_1024_1_IN_100 => FROM_STATE_REG_100 ,
										MUX_1024_1_IN_101 => FROM_STATE_REG_101 ,
										MUX_1024_1_IN_102 => FROM_STATE_REG_102 ,
										MUX_1024_1_IN_103 => FROM_STATE_REG_103 ,
										MUX_1024_1_IN_104 => FROM_STATE_REG_104 ,
										MUX_1024_1_IN_105 => FROM_STATE_REG_105 ,
										MUX_1024_1_IN_106 => FROM_STATE_REG_106 ,
										MUX_1024_1_IN_107 => FROM_STATE_REG_107 ,
										MUX_1024_1_IN_108 => FROM_STATE_REG_108 ,
										MUX_1024_1_IN_109 => FROM_STATE_REG_109 ,
										MUX_1024_1_IN_110 => FROM_STATE_REG_110 ,
										MUX_1024_1_IN_111 => FROM_STATE_REG_111 ,
										MUX_1024_1_IN_112 => FROM_STATE_REG_112 ,
										MUX_1024_1_IN_113 => FROM_STATE_REG_113 ,
										MUX_1024_1_IN_114 => FROM_STATE_REG_114 ,
										MUX_1024_1_IN_115 => FROM_STATE_REG_115 ,
										MUX_1024_1_IN_116 => FROM_STATE_REG_116 ,
										MUX_1024_1_IN_117 => FROM_STATE_REG_117 ,
										MUX_1024_1_IN_118 => FROM_STATE_REG_118 ,
										MUX_1024_1_IN_119 => FROM_STATE_REG_119 ,
										MUX_1024_1_IN_120 => FROM_STATE_REG_120 ,
										MUX_1024_1_IN_121 => FROM_STATE_REG_121 ,
										MUX_1024_1_IN_122 => FROM_STATE_REG_122 ,
										MUX_1024_1_IN_123 => FROM_STATE_REG_123 ,
										MUX_1024_1_IN_124 => FROM_STATE_REG_124 ,
										MUX_1024_1_IN_125 => FROM_STATE_REG_125 ,
										MUX_1024_1_IN_126 => FROM_STATE_REG_126 ,
										MUX_1024_1_IN_127 => FROM_STATE_REG_127 ,
										MUX_1024_1_IN_128 => FROM_STATE_REG_128 ,
										MUX_1024_1_IN_129 => FROM_STATE_REG_129 ,
										MUX_1024_1_IN_130 => FROM_STATE_REG_130 ,
										MUX_1024_1_IN_131 => FROM_STATE_REG_131 ,
										MUX_1024_1_IN_132 => FROM_STATE_REG_132 ,
										MUX_1024_1_IN_133 => FROM_STATE_REG_133 ,
										MUX_1024_1_IN_134 => FROM_STATE_REG_134 ,
										MUX_1024_1_IN_135 => FROM_STATE_REG_135 ,
										MUX_1024_1_IN_136 => FROM_STATE_REG_136 ,
										MUX_1024_1_IN_137 => FROM_STATE_REG_137 ,
										MUX_1024_1_IN_138 => FROM_STATE_REG_138 ,
										MUX_1024_1_IN_139 => FROM_STATE_REG_139 ,
										MUX_1024_1_IN_140 => FROM_STATE_REG_140 ,
										MUX_1024_1_IN_141 => FROM_STATE_REG_141 ,
										MUX_1024_1_IN_142 => FROM_STATE_REG_142 ,
										MUX_1024_1_IN_143 => FROM_STATE_REG_143 ,
										MUX_1024_1_IN_144 => FROM_STATE_REG_144 ,
										MUX_1024_1_IN_145 => FROM_STATE_REG_145 ,
										MUX_1024_1_IN_146 => FROM_STATE_REG_146 ,
										MUX_1024_1_IN_147 => FROM_STATE_REG_147 ,
										MUX_1024_1_IN_148 => FROM_STATE_REG_148 ,
										MUX_1024_1_IN_149 => FROM_STATE_REG_149 ,
										MUX_1024_1_IN_150 => FROM_STATE_REG_150 ,
										MUX_1024_1_IN_151 => FROM_STATE_REG_151 ,
										MUX_1024_1_IN_152 => FROM_STATE_REG_152 ,
										MUX_1024_1_IN_153 => FROM_STATE_REG_153 ,
										MUX_1024_1_IN_154 => FROM_STATE_REG_154 ,
										MUX_1024_1_IN_155 => FROM_STATE_REG_155 ,
										MUX_1024_1_IN_156 => FROM_STATE_REG_156 ,
										MUX_1024_1_IN_157 => FROM_STATE_REG_157 ,
										MUX_1024_1_IN_158 => FROM_STATE_REG_158 ,
										MUX_1024_1_IN_159 => FROM_STATE_REG_159 ,
										MUX_1024_1_IN_160 => FROM_STATE_REG_160 ,
										MUX_1024_1_IN_161 => FROM_STATE_REG_161 ,
										MUX_1024_1_IN_162 => FROM_STATE_REG_162 ,
										MUX_1024_1_IN_163 => FROM_STATE_REG_163 ,
										MUX_1024_1_IN_164 => FROM_STATE_REG_164 ,
										MUX_1024_1_IN_165 => FROM_STATE_REG_165 ,
										MUX_1024_1_IN_166 => FROM_STATE_REG_166 ,
										MUX_1024_1_IN_167 => FROM_STATE_REG_167 ,
										MUX_1024_1_IN_168 => FROM_STATE_REG_168 ,
										MUX_1024_1_IN_169 => FROM_STATE_REG_169 ,
										MUX_1024_1_IN_170 => FROM_STATE_REG_170 ,
										MUX_1024_1_IN_171 => FROM_STATE_REG_171 ,
										MUX_1024_1_IN_172 => FROM_STATE_REG_172 ,
										MUX_1024_1_IN_173 => FROM_STATE_REG_173 ,
										MUX_1024_1_IN_174 => FROM_STATE_REG_174 ,
										MUX_1024_1_IN_175 => FROM_STATE_REG_175 ,
										MUX_1024_1_IN_176 => FROM_STATE_REG_176 ,
										MUX_1024_1_IN_177 => FROM_STATE_REG_177 ,
										MUX_1024_1_IN_178 => FROM_STATE_REG_178 ,
										MUX_1024_1_IN_179 => FROM_STATE_REG_179 ,
										MUX_1024_1_IN_180 => FROM_STATE_REG_180 ,
										MUX_1024_1_IN_181 => FROM_STATE_REG_181 ,
										MUX_1024_1_IN_182 => FROM_STATE_REG_182 ,
										MUX_1024_1_IN_183 => FROM_STATE_REG_183 ,
										MUX_1024_1_IN_184 => FROM_STATE_REG_184 ,
										MUX_1024_1_IN_185 => FROM_STATE_REG_185 ,
										MUX_1024_1_IN_186 => FROM_STATE_REG_186 ,
										MUX_1024_1_IN_187 => FROM_STATE_REG_187 ,
										MUX_1024_1_IN_188 => FROM_STATE_REG_188 ,
										MUX_1024_1_IN_189 => FROM_STATE_REG_189 ,
										MUX_1024_1_IN_190 => FROM_STATE_REG_190 ,
										MUX_1024_1_IN_191 => FROM_STATE_REG_191 ,
										MUX_1024_1_IN_192 => FROM_STATE_REG_192 ,
										MUX_1024_1_IN_193 => FROM_STATE_REG_193 ,
										MUX_1024_1_IN_194 => FROM_STATE_REG_194 ,
										MUX_1024_1_IN_195 => FROM_STATE_REG_195 ,
										MUX_1024_1_IN_196 => FROM_STATE_REG_196 ,
										MUX_1024_1_IN_197 => FROM_STATE_REG_197 ,
										MUX_1024_1_IN_198 => FROM_STATE_REG_198 ,
										MUX_1024_1_IN_199 => FROM_STATE_REG_199 ,
										MUX_1024_1_IN_200 => FROM_STATE_REG_200 ,
										MUX_1024_1_IN_201 => FROM_STATE_REG_201 ,
										MUX_1024_1_IN_202 => FROM_STATE_REG_202 ,
										MUX_1024_1_IN_203 => FROM_STATE_REG_203 ,
										MUX_1024_1_IN_204 => FROM_STATE_REG_204 ,
										MUX_1024_1_IN_205 => FROM_STATE_REG_205 ,
										MUX_1024_1_IN_206 => FROM_STATE_REG_206 ,
										MUX_1024_1_IN_207 => FROM_STATE_REG_207 ,
										MUX_1024_1_IN_208 => FROM_STATE_REG_208 ,
										MUX_1024_1_IN_209 => FROM_STATE_REG_209 ,
										MUX_1024_1_IN_210 => FROM_STATE_REG_210 ,
										MUX_1024_1_IN_211 => FROM_STATE_REG_211 ,
										MUX_1024_1_IN_212 => FROM_STATE_REG_212 ,
										MUX_1024_1_IN_213 => FROM_STATE_REG_213 ,
										MUX_1024_1_IN_214 => FROM_STATE_REG_214 ,
										MUX_1024_1_IN_215 => FROM_STATE_REG_215 ,
										MUX_1024_1_IN_216 => FROM_STATE_REG_216 ,
										MUX_1024_1_IN_217 => FROM_STATE_REG_217 ,
										MUX_1024_1_IN_218 => FROM_STATE_REG_218 ,
										MUX_1024_1_IN_219 => FROM_STATE_REG_219 ,
										MUX_1024_1_IN_220 => FROM_STATE_REG_220 ,
										MUX_1024_1_IN_221 => FROM_STATE_REG_221 ,
										MUX_1024_1_IN_222 => FROM_STATE_REG_222 ,
										MUX_1024_1_IN_223 => FROM_STATE_REG_223 ,
										MUX_1024_1_IN_224 => FROM_STATE_REG_224 ,
										MUX_1024_1_IN_225 => FROM_STATE_REG_225 ,
										MUX_1024_1_IN_226 => FROM_STATE_REG_226 ,
										MUX_1024_1_IN_227 => FROM_STATE_REG_227 ,
										MUX_1024_1_IN_228 => FROM_STATE_REG_228 ,
										MUX_1024_1_IN_229 => FROM_STATE_REG_229 ,
										MUX_1024_1_IN_230 => FROM_STATE_REG_230 ,
										MUX_1024_1_IN_231 => FROM_STATE_REG_231 ,
										MUX_1024_1_IN_232 => FROM_STATE_REG_232 ,
										MUX_1024_1_IN_233 => FROM_STATE_REG_233 ,
										MUX_1024_1_IN_234 => FROM_STATE_REG_234 ,
										MUX_1024_1_IN_235 => FROM_STATE_REG_235 ,
										MUX_1024_1_IN_236 => FROM_STATE_REG_236 ,
										MUX_1024_1_IN_237 => FROM_STATE_REG_237 ,
										MUX_1024_1_IN_238 => FROM_STATE_REG_238 ,
										MUX_1024_1_IN_239 => FROM_STATE_REG_239 ,
										MUX_1024_1_IN_240 => FROM_STATE_REG_240 ,
										MUX_1024_1_IN_241 => FROM_STATE_REG_241 ,
										MUX_1024_1_IN_242 => FROM_STATE_REG_242 ,
										MUX_1024_1_IN_243 => FROM_STATE_REG_243 ,
										MUX_1024_1_IN_244 => FROM_STATE_REG_244 ,
										MUX_1024_1_IN_245 => FROM_STATE_REG_245 ,
										MUX_1024_1_IN_246 => FROM_STATE_REG_246 ,
										MUX_1024_1_IN_247 => FROM_STATE_REG_247 ,
										MUX_1024_1_IN_248 => FROM_STATE_REG_248 ,
										MUX_1024_1_IN_249 => FROM_STATE_REG_249 ,
										MUX_1024_1_IN_250 => FROM_STATE_REG_250 ,
										MUX_1024_1_IN_251 => FROM_STATE_REG_251 ,
										MUX_1024_1_IN_252 => FROM_STATE_REG_252 ,
										MUX_1024_1_IN_253 => FROM_STATE_REG_253 ,
										MUX_1024_1_IN_254 => FROM_STATE_REG_254 ,
										MUX_1024_1_IN_255 => FROM_STATE_REG_255 ,
										MUX_1024_1_IN_256 => FROM_STATE_REG_256 ,
										MUX_1024_1_IN_257 => FROM_STATE_REG_257 ,
										MUX_1024_1_IN_258 => FROM_STATE_REG_258 ,
										MUX_1024_1_IN_259 => FROM_STATE_REG_259 ,
										MUX_1024_1_IN_260 => FROM_STATE_REG_260 ,
										MUX_1024_1_IN_261 => FROM_STATE_REG_261 ,
										MUX_1024_1_IN_262 => FROM_STATE_REG_262 ,
										MUX_1024_1_IN_263 => FROM_STATE_REG_263 ,
										MUX_1024_1_IN_264 => FROM_STATE_REG_264 ,
										MUX_1024_1_IN_265 => FROM_STATE_REG_265 ,
										MUX_1024_1_IN_266 => FROM_STATE_REG_266 ,
										MUX_1024_1_IN_267 => FROM_STATE_REG_267 ,
										MUX_1024_1_IN_268 => FROM_STATE_REG_268 ,
										MUX_1024_1_IN_269 => FROM_STATE_REG_269 ,
										MUX_1024_1_IN_270 => FROM_STATE_REG_270 ,
										MUX_1024_1_IN_271 => FROM_STATE_REG_271 ,
										MUX_1024_1_IN_272 => FROM_STATE_REG_272 ,
										MUX_1024_1_IN_273 => FROM_STATE_REG_273 ,
										MUX_1024_1_IN_274 => FROM_STATE_REG_274 ,
										MUX_1024_1_IN_275 => FROM_STATE_REG_275 ,
										MUX_1024_1_IN_276 => FROM_STATE_REG_276 ,
										MUX_1024_1_IN_277 => FROM_STATE_REG_277 ,
										MUX_1024_1_IN_278 => FROM_STATE_REG_278 ,
										MUX_1024_1_IN_279 => FROM_STATE_REG_279 ,
										MUX_1024_1_IN_280 => FROM_STATE_REG_280 ,
										MUX_1024_1_IN_281 => FROM_STATE_REG_281 ,
										MUX_1024_1_IN_282 => FROM_STATE_REG_282 ,
										MUX_1024_1_IN_283 => FROM_STATE_REG_283 ,
										MUX_1024_1_IN_284 => FROM_STATE_REG_284 ,
										MUX_1024_1_IN_285 => FROM_STATE_REG_285 ,
										MUX_1024_1_IN_286 => FROM_STATE_REG_286 ,
										MUX_1024_1_IN_287 => FROM_STATE_REG_287 ,
										MUX_1024_1_IN_288 => FROM_STATE_REG_288 ,
										MUX_1024_1_IN_289 => FROM_STATE_REG_289 ,
										MUX_1024_1_IN_290 => FROM_STATE_REG_290 ,
										MUX_1024_1_IN_291 => FROM_STATE_REG_291 ,
										MUX_1024_1_IN_292 => FROM_STATE_REG_292 ,
										MUX_1024_1_IN_293 => FROM_STATE_REG_293 ,
										MUX_1024_1_IN_294 => FROM_STATE_REG_294 ,
										MUX_1024_1_IN_295 => FROM_STATE_REG_295 ,
										MUX_1024_1_IN_296 => FROM_STATE_REG_296 ,
										MUX_1024_1_IN_297 => FROM_STATE_REG_297 ,
										MUX_1024_1_IN_298 => FROM_STATE_REG_298 ,
										MUX_1024_1_IN_299 => FROM_STATE_REG_299 ,
										MUX_1024_1_IN_300 => FROM_STATE_REG_300 ,
										MUX_1024_1_IN_301 => FROM_STATE_REG_301 ,
										MUX_1024_1_IN_302 => FROM_STATE_REG_302 ,
										MUX_1024_1_IN_303 => FROM_STATE_REG_303 ,
										MUX_1024_1_IN_304 => FROM_STATE_REG_304 ,
										MUX_1024_1_IN_305 => FROM_STATE_REG_305 ,
										MUX_1024_1_IN_306 => FROM_STATE_REG_306 ,
										MUX_1024_1_IN_307 => FROM_STATE_REG_307 ,
										MUX_1024_1_IN_308 => FROM_STATE_REG_308 ,
										MUX_1024_1_IN_309 => FROM_STATE_REG_309 ,
										MUX_1024_1_IN_310 => FROM_STATE_REG_310 ,
										MUX_1024_1_IN_311 => FROM_STATE_REG_311 ,
										MUX_1024_1_IN_312 => FROM_STATE_REG_312 ,
										MUX_1024_1_IN_313 => FROM_STATE_REG_313 ,
										MUX_1024_1_IN_314 => FROM_STATE_REG_314 ,
										MUX_1024_1_IN_315 => FROM_STATE_REG_315 ,
										MUX_1024_1_IN_316 => FROM_STATE_REG_316 ,
										MUX_1024_1_IN_317 => FROM_STATE_REG_317 ,
										MUX_1024_1_IN_318 => FROM_STATE_REG_318 ,
										MUX_1024_1_IN_319 => FROM_STATE_REG_319 ,
										MUX_1024_1_IN_320 => FROM_STATE_REG_320 ,
										MUX_1024_1_IN_321 => FROM_STATE_REG_321 ,
										MUX_1024_1_IN_322 => FROM_STATE_REG_322 ,
										MUX_1024_1_IN_323 => FROM_STATE_REG_323 ,
										MUX_1024_1_IN_324 => FROM_STATE_REG_324 ,
										MUX_1024_1_IN_325 => FROM_STATE_REG_325 ,
										MUX_1024_1_IN_326 => FROM_STATE_REG_326 ,
										MUX_1024_1_IN_327 => FROM_STATE_REG_327 ,
										MUX_1024_1_IN_328 => FROM_STATE_REG_328 ,
										MUX_1024_1_IN_329 => FROM_STATE_REG_329 ,
										MUX_1024_1_IN_330 => FROM_STATE_REG_330 ,
										MUX_1024_1_IN_331 => FROM_STATE_REG_331 ,
										MUX_1024_1_IN_332 => FROM_STATE_REG_332 ,
										MUX_1024_1_IN_333 => FROM_STATE_REG_333 ,
										MUX_1024_1_IN_334 => FROM_STATE_REG_334 ,
										MUX_1024_1_IN_335 => FROM_STATE_REG_335 ,
										MUX_1024_1_IN_336 => FROM_STATE_REG_336 ,
										MUX_1024_1_IN_337 => FROM_STATE_REG_337 ,
										MUX_1024_1_IN_338 => FROM_STATE_REG_338 ,
										MUX_1024_1_IN_339 => FROM_STATE_REG_339 ,
										MUX_1024_1_IN_340 => FROM_STATE_REG_340 ,
										MUX_1024_1_IN_341 => FROM_STATE_REG_341 ,
										MUX_1024_1_IN_342 => FROM_STATE_REG_342 ,
										MUX_1024_1_IN_343 => FROM_STATE_REG_343 ,
										MUX_1024_1_IN_344 => FROM_STATE_REG_344 ,
										MUX_1024_1_IN_345 => FROM_STATE_REG_345 ,
										MUX_1024_1_IN_346 => FROM_STATE_REG_346 ,
										MUX_1024_1_IN_347 => FROM_STATE_REG_347 ,
										MUX_1024_1_IN_348 => FROM_STATE_REG_348 ,
										MUX_1024_1_IN_349 => FROM_STATE_REG_349 ,
										MUX_1024_1_IN_350 => FROM_STATE_REG_350 ,
										MUX_1024_1_IN_351 => FROM_STATE_REG_351 ,
										MUX_1024_1_IN_352 => FROM_STATE_REG_352 ,
										MUX_1024_1_IN_353 => FROM_STATE_REG_353 ,
										MUX_1024_1_IN_354 => FROM_STATE_REG_354 ,
										MUX_1024_1_IN_355 => FROM_STATE_REG_355 ,
										MUX_1024_1_IN_356 => FROM_STATE_REG_356 ,
										MUX_1024_1_IN_357 => FROM_STATE_REG_357 ,
										MUX_1024_1_IN_358 => FROM_STATE_REG_358 ,
										MUX_1024_1_IN_359 => FROM_STATE_REG_359 ,
										MUX_1024_1_IN_360 => FROM_STATE_REG_360 ,
										MUX_1024_1_IN_361 => FROM_STATE_REG_361 ,
										MUX_1024_1_IN_362 => FROM_STATE_REG_362 ,
										MUX_1024_1_IN_363 => FROM_STATE_REG_363 ,
										MUX_1024_1_IN_364 => FROM_STATE_REG_364 ,
										MUX_1024_1_IN_365 => FROM_STATE_REG_365 ,
										MUX_1024_1_IN_366 => FROM_STATE_REG_366 ,
										MUX_1024_1_IN_367 => FROM_STATE_REG_367 ,
										MUX_1024_1_IN_368 => FROM_STATE_REG_368 ,
										MUX_1024_1_IN_369 => FROM_STATE_REG_369 ,
										MUX_1024_1_IN_370 => FROM_STATE_REG_370 ,
										MUX_1024_1_IN_371 => FROM_STATE_REG_371 ,
										MUX_1024_1_IN_372 => FROM_STATE_REG_372 ,
										MUX_1024_1_IN_373 => FROM_STATE_REG_373 ,
										MUX_1024_1_IN_374 => FROM_STATE_REG_374 ,
										MUX_1024_1_IN_375 => FROM_STATE_REG_375 ,
										MUX_1024_1_IN_376 => FROM_STATE_REG_376 ,
										MUX_1024_1_IN_377 => FROM_STATE_REG_377 ,
										MUX_1024_1_IN_378 => FROM_STATE_REG_378 ,
										MUX_1024_1_IN_379 => FROM_STATE_REG_379 ,
										MUX_1024_1_IN_380 => FROM_STATE_REG_380 ,
										MUX_1024_1_IN_381 => FROM_STATE_REG_381 ,
										MUX_1024_1_IN_382 => FROM_STATE_REG_382 ,
										MUX_1024_1_IN_383 => FROM_STATE_REG_383 ,
										MUX_1024_1_IN_384 => FROM_STATE_REG_384 ,
										MUX_1024_1_IN_385 => FROM_STATE_REG_385 ,
										MUX_1024_1_IN_386 => FROM_STATE_REG_386 ,
										MUX_1024_1_IN_387 => FROM_STATE_REG_387 ,
										MUX_1024_1_IN_388 => FROM_STATE_REG_388 ,
										MUX_1024_1_IN_389 => FROM_STATE_REG_389 ,
										MUX_1024_1_IN_390 => FROM_STATE_REG_390 ,
										MUX_1024_1_IN_391 => FROM_STATE_REG_391 ,
										MUX_1024_1_IN_392 => FROM_STATE_REG_392 ,
										MUX_1024_1_IN_393 => FROM_STATE_REG_393 ,
										MUX_1024_1_IN_394 => FROM_STATE_REG_394 ,
										MUX_1024_1_IN_395 => FROM_STATE_REG_395 ,
										MUX_1024_1_IN_396 => FROM_STATE_REG_396 ,
										MUX_1024_1_IN_397 => FROM_STATE_REG_397 ,
										MUX_1024_1_IN_398 => FROM_STATE_REG_398 ,
										MUX_1024_1_IN_399 => FROM_STATE_REG_399 ,
										MUX_1024_1_IN_400 => FROM_STATE_REG_400 ,
										MUX_1024_1_IN_401 => FROM_STATE_REG_401 ,
										MUX_1024_1_IN_402 => FROM_STATE_REG_402 ,
										MUX_1024_1_IN_403 => FROM_STATE_REG_403 ,
										MUX_1024_1_IN_404 => FROM_STATE_REG_404 ,
										MUX_1024_1_IN_405 => FROM_STATE_REG_405 ,
										MUX_1024_1_IN_406 => FROM_STATE_REG_406 ,
										MUX_1024_1_IN_407 => FROM_STATE_REG_407 ,
										MUX_1024_1_IN_408 => FROM_STATE_REG_408 ,
										MUX_1024_1_IN_409 => FROM_STATE_REG_409 ,
										MUX_1024_1_IN_410 => FROM_STATE_REG_410 ,
										MUX_1024_1_IN_411 => FROM_STATE_REG_411 ,
										MUX_1024_1_IN_412 => FROM_STATE_REG_412 ,
										MUX_1024_1_IN_413 => FROM_STATE_REG_413 ,
										MUX_1024_1_IN_414 => FROM_STATE_REG_414 ,
										MUX_1024_1_IN_415 => FROM_STATE_REG_415 ,
										MUX_1024_1_IN_416 => FROM_STATE_REG_416 ,
										MUX_1024_1_IN_417 => FROM_STATE_REG_417 ,
										MUX_1024_1_IN_418 => FROM_STATE_REG_418 ,
										MUX_1024_1_IN_419 => FROM_STATE_REG_419 ,
										MUX_1024_1_IN_420 => FROM_STATE_REG_420 ,
										MUX_1024_1_IN_421 => FROM_STATE_REG_421 ,
										MUX_1024_1_IN_422 => FROM_STATE_REG_422 ,
										MUX_1024_1_IN_423 => FROM_STATE_REG_423 ,
										MUX_1024_1_IN_424 => FROM_STATE_REG_424 ,
										MUX_1024_1_IN_425 => FROM_STATE_REG_425 ,
										MUX_1024_1_IN_426 => FROM_STATE_REG_426 ,
										MUX_1024_1_IN_427 => FROM_STATE_REG_427 ,
										MUX_1024_1_IN_428 => FROM_STATE_REG_428 ,
										MUX_1024_1_IN_429 => FROM_STATE_REG_429 ,
										MUX_1024_1_IN_430 => FROM_STATE_REG_430 ,
										MUX_1024_1_IN_431 => FROM_STATE_REG_431 ,
										MUX_1024_1_IN_432 => FROM_STATE_REG_432 ,
										MUX_1024_1_IN_433 => FROM_STATE_REG_433 ,
										MUX_1024_1_IN_434 => FROM_STATE_REG_434 ,
										MUX_1024_1_IN_435 => FROM_STATE_REG_435 ,
										MUX_1024_1_IN_436 => FROM_STATE_REG_436 ,
										MUX_1024_1_IN_437 => FROM_STATE_REG_437 ,
										MUX_1024_1_IN_438 => FROM_STATE_REG_438 ,
										MUX_1024_1_IN_439 => FROM_STATE_REG_439 ,
										MUX_1024_1_IN_440 => FROM_STATE_REG_440 ,
										MUX_1024_1_IN_441 => FROM_STATE_REG_441 ,
										MUX_1024_1_IN_442 => FROM_STATE_REG_442 ,
										MUX_1024_1_IN_443 => FROM_STATE_REG_443 ,
										MUX_1024_1_IN_444 => FROM_STATE_REG_444 ,
										MUX_1024_1_IN_445 => FROM_STATE_REG_445 ,
										MUX_1024_1_IN_446 => FROM_STATE_REG_446 ,
										MUX_1024_1_IN_447 => FROM_STATE_REG_447 ,
										MUX_1024_1_IN_448 => FROM_STATE_REG_448 ,
										MUX_1024_1_IN_449 => FROM_STATE_REG_449 ,
										MUX_1024_1_IN_450 => FROM_STATE_REG_450 ,
										MUX_1024_1_IN_451 => FROM_STATE_REG_451 ,
										MUX_1024_1_IN_452 => FROM_STATE_REG_452 ,
										MUX_1024_1_IN_453 => FROM_STATE_REG_453 ,
										MUX_1024_1_IN_454 => FROM_STATE_REG_454 ,
										MUX_1024_1_IN_455 => FROM_STATE_REG_455 ,
										MUX_1024_1_IN_456 => FROM_STATE_REG_456 ,
										MUX_1024_1_IN_457 => FROM_STATE_REG_457 ,
										MUX_1024_1_IN_458 => FROM_STATE_REG_458 ,
										MUX_1024_1_IN_459 => FROM_STATE_REG_459 ,
										MUX_1024_1_IN_460 => FROM_STATE_REG_460 ,
										MUX_1024_1_IN_461 => FROM_STATE_REG_461 ,
										MUX_1024_1_IN_462 => FROM_STATE_REG_462 ,
										MUX_1024_1_IN_463 => FROM_STATE_REG_463 ,
										MUX_1024_1_IN_464 => FROM_STATE_REG_464 ,
										MUX_1024_1_IN_465 => FROM_STATE_REG_465 ,
										MUX_1024_1_IN_466 => FROM_STATE_REG_466 ,
										MUX_1024_1_IN_467 => FROM_STATE_REG_467 ,
										MUX_1024_1_IN_468 => FROM_STATE_REG_468 ,
										MUX_1024_1_IN_469 => FROM_STATE_REG_469 ,
										MUX_1024_1_IN_470 => FROM_STATE_REG_470 ,
										MUX_1024_1_IN_471 => FROM_STATE_REG_471 ,
										MUX_1024_1_IN_472 => FROM_STATE_REG_472 ,
										MUX_1024_1_IN_473 => FROM_STATE_REG_473 ,
										MUX_1024_1_IN_474 => FROM_STATE_REG_474 ,
										MUX_1024_1_IN_475 => FROM_STATE_REG_475 ,
										MUX_1024_1_IN_476 => FROM_STATE_REG_476 ,
										MUX_1024_1_IN_477 => FROM_STATE_REG_477 ,
										MUX_1024_1_IN_478 => FROM_STATE_REG_478 ,
										MUX_1024_1_IN_479 => FROM_STATE_REG_479 ,
										MUX_1024_1_IN_480 => FROM_STATE_REG_480 ,
										MUX_1024_1_IN_481 => FROM_STATE_REG_481 ,
										MUX_1024_1_IN_482 => FROM_STATE_REG_482 ,
										MUX_1024_1_IN_483 => FROM_STATE_REG_483 ,
										MUX_1024_1_IN_484 => FROM_STATE_REG_484 ,
										MUX_1024_1_IN_485 => FROM_STATE_REG_485 ,
										MUX_1024_1_IN_486 => FROM_STATE_REG_486 ,
										MUX_1024_1_IN_487 => FROM_STATE_REG_487 ,
										MUX_1024_1_IN_488 => FROM_STATE_REG_488 ,
										MUX_1024_1_IN_489 => FROM_STATE_REG_489 ,
										MUX_1024_1_IN_490 => FROM_STATE_REG_490 ,
										MUX_1024_1_IN_491 => FROM_STATE_REG_491 ,
										MUX_1024_1_IN_492 => FROM_STATE_REG_492 ,
										MUX_1024_1_IN_493 => FROM_STATE_REG_493 ,
										MUX_1024_1_IN_494 => FROM_STATE_REG_494 ,
										MUX_1024_1_IN_495 => FROM_STATE_REG_495 ,
										MUX_1024_1_IN_496 => FROM_STATE_REG_496 ,
										MUX_1024_1_IN_497 => FROM_STATE_REG_497 ,
										MUX_1024_1_IN_498 => FROM_STATE_REG_498 ,
										MUX_1024_1_IN_499 => FROM_STATE_REG_499 ,
										MUX_1024_1_IN_500 => FROM_STATE_REG_500 ,
										MUX_1024_1_IN_501 => FROM_STATE_REG_501 ,
										MUX_1024_1_IN_502 => FROM_STATE_REG_502 ,
										MUX_1024_1_IN_503 => FROM_STATE_REG_503 ,
										MUX_1024_1_IN_504 => FROM_STATE_REG_504 ,
										MUX_1024_1_IN_505 => FROM_STATE_REG_505 ,
										MUX_1024_1_IN_506 => FROM_STATE_REG_506 ,
										MUX_1024_1_IN_507 => FROM_STATE_REG_507 ,
										MUX_1024_1_IN_508 => FROM_STATE_REG_508 ,
										MUX_1024_1_IN_509 => FROM_STATE_REG_509 ,
										MUX_1024_1_IN_510 => FROM_STATE_REG_510 ,
										MUX_1024_1_IN_511 => FROM_STATE_REG_511 ,
										MUX_1024_1_IN_512 => FROM_STATE_REG_512 ,
										MUX_1024_1_IN_513 => FROM_STATE_REG_513 ,
										MUX_1024_1_IN_514 => FROM_STATE_REG_514 ,
										MUX_1024_1_IN_515 => FROM_STATE_REG_515 ,
										MUX_1024_1_IN_516 => FROM_STATE_REG_516 ,
										MUX_1024_1_IN_517 => FROM_STATE_REG_517 ,
										MUX_1024_1_IN_518 => FROM_STATE_REG_518 ,
										MUX_1024_1_IN_519 => FROM_STATE_REG_519 ,
										MUX_1024_1_IN_520 => FROM_STATE_REG_520 ,
										MUX_1024_1_IN_521 => FROM_STATE_REG_521 ,
										MUX_1024_1_IN_522 => FROM_STATE_REG_522 ,
										MUX_1024_1_IN_523 => FROM_STATE_REG_523 ,
										MUX_1024_1_IN_524 => FROM_STATE_REG_524 ,
										MUX_1024_1_IN_525 => FROM_STATE_REG_525 ,
										MUX_1024_1_IN_526 => FROM_STATE_REG_526 ,
										MUX_1024_1_IN_527 => FROM_STATE_REG_527 ,
										MUX_1024_1_IN_528 => FROM_STATE_REG_528 ,
										MUX_1024_1_IN_529 => FROM_STATE_REG_529 ,
										MUX_1024_1_IN_530 => FROM_STATE_REG_530 ,
										MUX_1024_1_IN_531 => FROM_STATE_REG_531 ,
										MUX_1024_1_IN_532 => FROM_STATE_REG_532 ,
										MUX_1024_1_IN_533 => FROM_STATE_REG_533 ,
										MUX_1024_1_IN_534 => FROM_STATE_REG_534 ,
										MUX_1024_1_IN_535 => FROM_STATE_REG_535 ,
										MUX_1024_1_IN_536 => FROM_STATE_REG_536 ,
										MUX_1024_1_IN_537 => FROM_STATE_REG_537 ,
										MUX_1024_1_IN_538 => FROM_STATE_REG_538 ,
										MUX_1024_1_IN_539 => FROM_STATE_REG_539 ,
										MUX_1024_1_IN_540 => FROM_STATE_REG_540 ,
										MUX_1024_1_IN_541 => FROM_STATE_REG_541 ,
										MUX_1024_1_IN_542 => FROM_STATE_REG_542 ,
										MUX_1024_1_IN_543 => FROM_STATE_REG_543 ,
										MUX_1024_1_IN_544 => FROM_STATE_REG_544 ,
										MUX_1024_1_IN_545 => FROM_STATE_REG_545 ,
										MUX_1024_1_IN_546 => FROM_STATE_REG_546 ,
										MUX_1024_1_IN_547 => FROM_STATE_REG_547 ,
										MUX_1024_1_IN_548 => FROM_STATE_REG_548 ,
										MUX_1024_1_IN_549 => FROM_STATE_REG_549 ,
										MUX_1024_1_IN_550 => FROM_STATE_REG_550 ,
										MUX_1024_1_IN_551 => FROM_STATE_REG_551 ,
										MUX_1024_1_IN_552 => FROM_STATE_REG_552 ,
										MUX_1024_1_IN_553 => FROM_STATE_REG_553 ,
										MUX_1024_1_IN_554 => FROM_STATE_REG_554 ,
										MUX_1024_1_IN_555 => FROM_STATE_REG_555 ,
										MUX_1024_1_IN_556 => FROM_STATE_REG_556 ,
										MUX_1024_1_IN_557 => FROM_STATE_REG_557 ,
										MUX_1024_1_IN_558 => FROM_STATE_REG_558 ,
										MUX_1024_1_IN_559 => FROM_STATE_REG_559 ,
										MUX_1024_1_IN_560 => FROM_STATE_REG_560 ,
										MUX_1024_1_IN_561 => FROM_STATE_REG_561 ,
										MUX_1024_1_IN_562 => FROM_STATE_REG_562 ,
										MUX_1024_1_IN_563 => FROM_STATE_REG_563 ,
										MUX_1024_1_IN_564 => FROM_STATE_REG_564 ,
										MUX_1024_1_IN_565 => FROM_STATE_REG_565 ,
										MUX_1024_1_IN_566 => FROM_STATE_REG_566 ,
										MUX_1024_1_IN_567 => FROM_STATE_REG_567 ,
										MUX_1024_1_IN_568 => FROM_STATE_REG_568 ,
										MUX_1024_1_IN_569 => FROM_STATE_REG_569 ,
										MUX_1024_1_IN_570 => FROM_STATE_REG_570 ,
										MUX_1024_1_IN_571 => FROM_STATE_REG_571 ,
										MUX_1024_1_IN_572 => FROM_STATE_REG_572 ,
										MUX_1024_1_IN_573 => FROM_STATE_REG_573 ,
										MUX_1024_1_IN_574 => FROM_STATE_REG_574 ,
										MUX_1024_1_IN_575 => FROM_STATE_REG_575 ,
										MUX_1024_1_IN_576 => FROM_STATE_REG_576 ,
										MUX_1024_1_IN_577 => FROM_STATE_REG_577 ,
										MUX_1024_1_IN_578 => FROM_STATE_REG_578 ,
										MUX_1024_1_IN_579 => FROM_STATE_REG_579 ,
										MUX_1024_1_IN_580 => FROM_STATE_REG_580 ,
										MUX_1024_1_IN_581 => FROM_STATE_REG_581 ,
										MUX_1024_1_IN_582 => FROM_STATE_REG_582 ,
										MUX_1024_1_IN_583 => FROM_STATE_REG_583 ,
										MUX_1024_1_IN_584 => FROM_STATE_REG_584 ,
										MUX_1024_1_IN_585 => FROM_STATE_REG_585 ,
										MUX_1024_1_IN_586 => FROM_STATE_REG_586 ,
										MUX_1024_1_IN_587 => FROM_STATE_REG_587 ,
										MUX_1024_1_IN_588 => FROM_STATE_REG_588 ,
										MUX_1024_1_IN_589 => FROM_STATE_REG_589 ,
										MUX_1024_1_IN_590 => FROM_STATE_REG_590 ,
										MUX_1024_1_IN_591 => FROM_STATE_REG_591 ,
										MUX_1024_1_IN_592 => FROM_STATE_REG_592 ,
										MUX_1024_1_IN_593 => FROM_STATE_REG_593 ,
										MUX_1024_1_IN_594 => FROM_STATE_REG_594 ,
										MUX_1024_1_IN_595 => FROM_STATE_REG_595 ,
										MUX_1024_1_IN_596 => FROM_STATE_REG_596 ,
										MUX_1024_1_IN_597 => FROM_STATE_REG_597 ,
										MUX_1024_1_IN_598 => FROM_STATE_REG_598 ,
										MUX_1024_1_IN_599 => FROM_STATE_REG_599 ,
										MUX_1024_1_IN_600 => FROM_STATE_REG_600 ,
										MUX_1024_1_IN_601 => FROM_STATE_REG_601 ,
										MUX_1024_1_IN_602 => FROM_STATE_REG_602 ,
										MUX_1024_1_IN_603 => FROM_STATE_REG_603 ,
										MUX_1024_1_IN_604 => FROM_STATE_REG_604 ,
										MUX_1024_1_IN_605 => FROM_STATE_REG_605 ,
										MUX_1024_1_IN_606 => FROM_STATE_REG_606 ,
										MUX_1024_1_IN_607 => FROM_STATE_REG_607 ,
										MUX_1024_1_IN_608 => FROM_STATE_REG_608 ,
										MUX_1024_1_IN_609 => FROM_STATE_REG_609 ,
										MUX_1024_1_IN_610 => FROM_STATE_REG_610 ,
										MUX_1024_1_IN_611 => FROM_STATE_REG_611 ,
										MUX_1024_1_IN_612 => FROM_STATE_REG_612 ,
										MUX_1024_1_IN_613 => FROM_STATE_REG_613 ,
										MUX_1024_1_IN_614 => FROM_STATE_REG_614 ,
										MUX_1024_1_IN_615 => FROM_STATE_REG_615 ,
										MUX_1024_1_IN_616 => FROM_STATE_REG_616 ,
										MUX_1024_1_IN_617 => FROM_STATE_REG_617 ,
										MUX_1024_1_IN_618 => FROM_STATE_REG_618 ,
										MUX_1024_1_IN_619 => FROM_STATE_REG_619 ,
										MUX_1024_1_IN_620 => FROM_STATE_REG_620 ,
										MUX_1024_1_IN_621 => FROM_STATE_REG_621 ,
										MUX_1024_1_IN_622 => FROM_STATE_REG_622 ,
										MUX_1024_1_IN_623 => FROM_STATE_REG_623 ,
										MUX_1024_1_IN_624 => FROM_STATE_REG_624 ,
										MUX_1024_1_IN_625 => FROM_STATE_REG_625 ,
										MUX_1024_1_IN_626 => FROM_STATE_REG_626 ,
										MUX_1024_1_IN_627 => FROM_STATE_REG_627 ,
										MUX_1024_1_IN_628 => FROM_STATE_REG_628 ,
										MUX_1024_1_IN_629 => FROM_STATE_REG_629 ,
										MUX_1024_1_IN_630 => FROM_STATE_REG_630 ,
										MUX_1024_1_IN_631 => FROM_STATE_REG_631 ,
										MUX_1024_1_IN_632 => FROM_STATE_REG_632 ,
										MUX_1024_1_IN_633 => FROM_STATE_REG_633 ,
										MUX_1024_1_IN_634 => FROM_STATE_REG_634 ,
										MUX_1024_1_IN_635 => FROM_STATE_REG_635 ,
										MUX_1024_1_IN_636 => FROM_STATE_REG_636 ,
										MUX_1024_1_IN_637 => FROM_STATE_REG_637 ,
										MUX_1024_1_IN_638 => FROM_STATE_REG_638 ,
										MUX_1024_1_IN_639 => FROM_STATE_REG_639 ,
										MUX_1024_1_IN_640 => FROM_STATE_REG_640 ,
										MUX_1024_1_IN_641 => FROM_STATE_REG_641 ,
										MUX_1024_1_IN_642 => FROM_STATE_REG_642 ,
										MUX_1024_1_IN_643 => FROM_STATE_REG_643 ,
										MUX_1024_1_IN_644 => FROM_STATE_REG_644 ,
										MUX_1024_1_IN_645 => FROM_STATE_REG_645 ,
										MUX_1024_1_IN_646 => FROM_STATE_REG_646 ,
										MUX_1024_1_IN_647 => FROM_STATE_REG_647 ,
										MUX_1024_1_IN_648 => FROM_STATE_REG_648 ,
										MUX_1024_1_IN_649 => FROM_STATE_REG_649 ,
										MUX_1024_1_IN_650 => FROM_STATE_REG_650 ,
										MUX_1024_1_IN_651 => FROM_STATE_REG_651 ,
										MUX_1024_1_IN_652 => FROM_STATE_REG_652 ,
										MUX_1024_1_IN_653 => FROM_STATE_REG_653 ,
										MUX_1024_1_IN_654 => FROM_STATE_REG_654 ,
										MUX_1024_1_IN_655 => FROM_STATE_REG_655 ,
										MUX_1024_1_IN_656 => FROM_STATE_REG_656 ,
										MUX_1024_1_IN_657 => FROM_STATE_REG_657 ,
										MUX_1024_1_IN_658 => FROM_STATE_REG_658 ,
										MUX_1024_1_IN_659 => FROM_STATE_REG_659 ,
										MUX_1024_1_IN_660 => FROM_STATE_REG_660 ,
										MUX_1024_1_IN_661 => FROM_STATE_REG_661 ,
										MUX_1024_1_IN_662 => FROM_STATE_REG_662 ,
										MUX_1024_1_IN_663 => FROM_STATE_REG_663 ,
										MUX_1024_1_IN_664 => FROM_STATE_REG_664 ,
										MUX_1024_1_IN_665 => FROM_STATE_REG_665 ,
										MUX_1024_1_IN_666 => FROM_STATE_REG_666 ,
										MUX_1024_1_IN_667 => FROM_STATE_REG_667 ,
										MUX_1024_1_IN_668 => FROM_STATE_REG_668 ,
										MUX_1024_1_IN_669 => FROM_STATE_REG_669 ,
										MUX_1024_1_IN_670 => FROM_STATE_REG_670 ,
										MUX_1024_1_IN_671 => FROM_STATE_REG_671 ,
										MUX_1024_1_IN_672 => FROM_STATE_REG_672 ,
										MUX_1024_1_IN_673 => FROM_STATE_REG_673 ,
										MUX_1024_1_IN_674 => FROM_STATE_REG_674 ,
										MUX_1024_1_IN_675 => FROM_STATE_REG_675 ,
										MUX_1024_1_IN_676 => FROM_STATE_REG_676 ,
										MUX_1024_1_IN_677 => FROM_STATE_REG_677 ,
										MUX_1024_1_IN_678 => FROM_STATE_REG_678 ,
										MUX_1024_1_IN_679 => FROM_STATE_REG_679 ,
										MUX_1024_1_IN_680 => FROM_STATE_REG_680 ,
										MUX_1024_1_IN_681 => FROM_STATE_REG_681 ,
										MUX_1024_1_IN_682 => FROM_STATE_REG_682 ,
										MUX_1024_1_IN_683 => FROM_STATE_REG_683 ,
										MUX_1024_1_IN_684 => FROM_STATE_REG_684 ,
										MUX_1024_1_IN_685 => FROM_STATE_REG_685 ,
										MUX_1024_1_IN_686 => FROM_STATE_REG_686 ,
										MUX_1024_1_IN_687 => FROM_STATE_REG_687 ,
										MUX_1024_1_IN_688 => FROM_STATE_REG_688 ,
										MUX_1024_1_IN_689 => FROM_STATE_REG_689 ,
										MUX_1024_1_IN_690 => FROM_STATE_REG_690 ,
										MUX_1024_1_IN_691 => FROM_STATE_REG_691 ,
										MUX_1024_1_IN_692 => FROM_STATE_REG_692 ,
										MUX_1024_1_IN_693 => FROM_STATE_REG_693 ,
										MUX_1024_1_IN_694 => FROM_STATE_REG_694 ,
										MUX_1024_1_IN_695 => FROM_STATE_REG_695 ,
										MUX_1024_1_IN_696 => FROM_STATE_REG_696 ,
										MUX_1024_1_IN_697 => FROM_STATE_REG_697 ,
										MUX_1024_1_IN_698 => FROM_STATE_REG_698 ,
										MUX_1024_1_IN_699 => FROM_STATE_REG_699 ,
										MUX_1024_1_IN_700 => FROM_STATE_REG_700 ,
										MUX_1024_1_IN_701 => FROM_STATE_REG_701 ,
										MUX_1024_1_IN_702 => FROM_STATE_REG_702 ,
										MUX_1024_1_IN_703 => FROM_STATE_REG_703 ,
										MUX_1024_1_IN_704 => FROM_STATE_REG_704 ,
										MUX_1024_1_IN_705 => FROM_STATE_REG_705 ,
										MUX_1024_1_IN_706 => FROM_STATE_REG_706 ,
										MUX_1024_1_IN_707 => FROM_STATE_REG_707 ,
										MUX_1024_1_IN_708 => FROM_STATE_REG_708 ,
										MUX_1024_1_IN_709 => FROM_STATE_REG_709 ,
										MUX_1024_1_IN_710 => FROM_STATE_REG_710 ,
										MUX_1024_1_IN_711 => FROM_STATE_REG_711 ,
										MUX_1024_1_IN_712 => FROM_STATE_REG_712 ,
										MUX_1024_1_IN_713 => FROM_STATE_REG_713 ,
										MUX_1024_1_IN_714 => FROM_STATE_REG_714 ,
										MUX_1024_1_IN_715 => FROM_STATE_REG_715 ,
										MUX_1024_1_IN_716 => FROM_STATE_REG_716 ,
										MUX_1024_1_IN_717 => FROM_STATE_REG_717 ,
										MUX_1024_1_IN_718 => FROM_STATE_REG_718 ,
										MUX_1024_1_IN_719 => FROM_STATE_REG_719 ,
										MUX_1024_1_IN_720 => FROM_STATE_REG_720 ,
										MUX_1024_1_IN_721 => FROM_STATE_REG_721 ,
										MUX_1024_1_IN_722 => FROM_STATE_REG_722 ,
										MUX_1024_1_IN_723 => FROM_STATE_REG_723 ,
										MUX_1024_1_IN_724 => FROM_STATE_REG_724 ,
										MUX_1024_1_IN_725 => FROM_STATE_REG_725 ,
										MUX_1024_1_IN_726 => FROM_STATE_REG_726 ,
										MUX_1024_1_IN_727 => FROM_STATE_REG_727 ,
										MUX_1024_1_IN_728 => FROM_STATE_REG_728 ,
										MUX_1024_1_IN_729 => FROM_STATE_REG_729 ,
										MUX_1024_1_IN_730 => FROM_STATE_REG_730 ,
										MUX_1024_1_IN_731 => FROM_STATE_REG_731 ,
										MUX_1024_1_IN_732 => FROM_STATE_REG_732 ,
										MUX_1024_1_IN_733 => FROM_STATE_REG_733 ,
										MUX_1024_1_IN_734 => FROM_STATE_REG_734 ,
										MUX_1024_1_IN_735 => FROM_STATE_REG_735 ,
										MUX_1024_1_IN_736 => FROM_STATE_REG_736 ,
										MUX_1024_1_IN_737 => FROM_STATE_REG_737 ,
										MUX_1024_1_IN_738 => FROM_STATE_REG_738 ,
										MUX_1024_1_IN_739 => FROM_STATE_REG_739 ,
										MUX_1024_1_IN_740 => FROM_STATE_REG_740 ,
										MUX_1024_1_IN_741 => FROM_STATE_REG_741 ,
										MUX_1024_1_IN_742 => FROM_STATE_REG_742 ,
										MUX_1024_1_IN_743 => FROM_STATE_REG_743 ,
										MUX_1024_1_IN_744 => FROM_STATE_REG_744 ,
										MUX_1024_1_IN_745 => FROM_STATE_REG_745 ,
										MUX_1024_1_IN_746 => FROM_STATE_REG_746 ,
										MUX_1024_1_IN_747 => FROM_STATE_REG_747 ,
										MUX_1024_1_IN_748 => FROM_STATE_REG_748 ,
										MUX_1024_1_IN_749 => FROM_STATE_REG_749 ,
										MUX_1024_1_IN_750 => FROM_STATE_REG_750 ,
										MUX_1024_1_IN_751 => FROM_STATE_REG_751 ,
										MUX_1024_1_IN_752 => FROM_STATE_REG_752 ,
										MUX_1024_1_IN_753 => FROM_STATE_REG_753 ,
										MUX_1024_1_IN_754 => FROM_STATE_REG_754 ,
										MUX_1024_1_IN_755 => FROM_STATE_REG_755 ,
										MUX_1024_1_IN_756 => FROM_STATE_REG_756 ,
										MUX_1024_1_IN_757 => FROM_STATE_REG_757 ,
										MUX_1024_1_IN_758 => FROM_STATE_REG_758 ,
										MUX_1024_1_IN_759 => FROM_STATE_REG_759 ,
										MUX_1024_1_IN_760 => FROM_STATE_REG_760 ,
										MUX_1024_1_IN_761 => FROM_STATE_REG_761 ,
										MUX_1024_1_IN_762 => FROM_STATE_REG_762 ,
										MUX_1024_1_IN_763 => FROM_STATE_REG_763 ,
										MUX_1024_1_IN_764 => FROM_STATE_REG_764 ,
										MUX_1024_1_IN_765 => FROM_STATE_REG_765 ,
										MUX_1024_1_IN_766 => FROM_STATE_REG_766 ,
										MUX_1024_1_IN_767 => FROM_STATE_REG_767 ,
										MUX_1024_1_IN_768 => FROM_STATE_REG_768 ,
										MUX_1024_1_IN_769 => FROM_STATE_REG_769 ,
										MUX_1024_1_IN_770 => FROM_STATE_REG_770 ,
										MUX_1024_1_IN_771 => FROM_STATE_REG_771 ,
										MUX_1024_1_IN_772 => FROM_STATE_REG_772 ,
										MUX_1024_1_IN_773 => FROM_STATE_REG_773 ,
										MUX_1024_1_IN_774 => FROM_STATE_REG_774 ,
										MUX_1024_1_IN_775 => FROM_STATE_REG_775 ,
										MUX_1024_1_IN_776 => FROM_STATE_REG_776 ,
										MUX_1024_1_IN_777 => FROM_STATE_REG_777 ,
										MUX_1024_1_IN_778 => FROM_STATE_REG_778 ,
										MUX_1024_1_IN_779 => FROM_STATE_REG_779 ,
										MUX_1024_1_IN_780 => FROM_STATE_REG_780 ,
										MUX_1024_1_IN_781 => FROM_STATE_REG_781 ,
										MUX_1024_1_IN_782 => FROM_STATE_REG_782 ,
										MUX_1024_1_IN_783 => FROM_STATE_REG_783 ,
										MUX_1024_1_IN_784 => FROM_STATE_REG_784 ,
										MUX_1024_1_IN_785 => FROM_STATE_REG_785 ,
										MUX_1024_1_IN_786 => FROM_STATE_REG_786 ,
										MUX_1024_1_IN_787 => FROM_STATE_REG_787 ,
										MUX_1024_1_IN_788 => FROM_STATE_REG_788 ,
										MUX_1024_1_IN_789 => FROM_STATE_REG_789 ,
										MUX_1024_1_IN_790 => FROM_STATE_REG_790 ,
										MUX_1024_1_IN_791 => FROM_STATE_REG_791 ,
										MUX_1024_1_IN_792 => FROM_STATE_REG_792 ,
										MUX_1024_1_IN_793 => FROM_STATE_REG_793 ,
										MUX_1024_1_IN_794 => FROM_STATE_REG_794 ,
										MUX_1024_1_IN_795 => FROM_STATE_REG_795 ,
										MUX_1024_1_IN_796 => FROM_STATE_REG_796 ,
										MUX_1024_1_IN_797 => FROM_STATE_REG_797 ,
										MUX_1024_1_IN_798 => FROM_STATE_REG_798 ,
										MUX_1024_1_IN_799 => FROM_STATE_REG_799 ,
										MUX_1024_1_IN_800 => FROM_STATE_REG_800 ,
										MUX_1024_1_IN_801 => FROM_STATE_REG_801 ,
										MUX_1024_1_IN_802 => FROM_STATE_REG_802 ,
										MUX_1024_1_IN_803 => FROM_STATE_REG_803 ,
										MUX_1024_1_IN_804 => FROM_STATE_REG_804 ,
										MUX_1024_1_IN_805 => FROM_STATE_REG_805 ,
										MUX_1024_1_IN_806 => FROM_STATE_REG_806 ,
										MUX_1024_1_IN_807 => FROM_STATE_REG_807 ,
										MUX_1024_1_IN_808 => FROM_STATE_REG_808 ,
										MUX_1024_1_IN_809 => FROM_STATE_REG_809 ,
										MUX_1024_1_IN_810 => FROM_STATE_REG_810 ,
										MUX_1024_1_IN_811 => FROM_STATE_REG_811 ,
										MUX_1024_1_IN_812 => FROM_STATE_REG_812 ,
										MUX_1024_1_IN_813 => FROM_STATE_REG_813 ,
										MUX_1024_1_IN_814 => FROM_STATE_REG_814 ,
										MUX_1024_1_IN_815 => FROM_STATE_REG_815 ,
										MUX_1024_1_IN_816 => FROM_STATE_REG_816 ,
										MUX_1024_1_IN_817 => FROM_STATE_REG_817 ,
										MUX_1024_1_IN_818 => FROM_STATE_REG_818 ,
										MUX_1024_1_IN_819 => FROM_STATE_REG_819 ,
										MUX_1024_1_IN_820 => FROM_STATE_REG_820 ,
										MUX_1024_1_IN_821 => FROM_STATE_REG_821 ,
										MUX_1024_1_IN_822 => FROM_STATE_REG_822 ,
										MUX_1024_1_IN_823 => FROM_STATE_REG_823 ,
										MUX_1024_1_IN_824 => FROM_STATE_REG_824 ,
										MUX_1024_1_IN_825 => FROM_STATE_REG_825 ,
										MUX_1024_1_IN_826 => FROM_STATE_REG_826 ,
										MUX_1024_1_IN_827 => FROM_STATE_REG_827 ,
										MUX_1024_1_IN_828 => FROM_STATE_REG_828 ,
										MUX_1024_1_IN_829 => FROM_STATE_REG_829 ,
										MUX_1024_1_IN_830 => FROM_STATE_REG_830 ,
										MUX_1024_1_IN_831 => FROM_STATE_REG_831 ,
										MUX_1024_1_IN_832 => FROM_STATE_REG_832 ,
										MUX_1024_1_IN_833 => FROM_STATE_REG_833 ,
										MUX_1024_1_IN_834 => FROM_STATE_REG_834 ,
										MUX_1024_1_IN_835 => FROM_STATE_REG_835 ,
										MUX_1024_1_IN_836 => FROM_STATE_REG_836 ,
										MUX_1024_1_IN_837 => FROM_STATE_REG_837 ,
										MUX_1024_1_IN_838 => FROM_STATE_REG_838 ,
										MUX_1024_1_IN_839 => FROM_STATE_REG_839 ,
										MUX_1024_1_IN_840 => FROM_STATE_REG_840 ,
										MUX_1024_1_IN_841 => FROM_STATE_REG_841 ,
										MUX_1024_1_IN_842 => FROM_STATE_REG_842 ,
										MUX_1024_1_IN_843 => FROM_STATE_REG_843 ,
										MUX_1024_1_IN_844 => FROM_STATE_REG_844 ,
										MUX_1024_1_IN_845 => FROM_STATE_REG_845 ,
										MUX_1024_1_IN_846 => FROM_STATE_REG_846 ,
										MUX_1024_1_IN_847 => FROM_STATE_REG_847 ,
										MUX_1024_1_IN_848 => FROM_STATE_REG_848 ,
										MUX_1024_1_IN_849 => FROM_STATE_REG_849 ,
										MUX_1024_1_IN_850 => FROM_STATE_REG_850 ,
										MUX_1024_1_IN_851 => FROM_STATE_REG_851 ,
										MUX_1024_1_IN_852 => FROM_STATE_REG_852 ,
										MUX_1024_1_IN_853 => FROM_STATE_REG_853 ,
										MUX_1024_1_IN_854 => FROM_STATE_REG_854 ,
										MUX_1024_1_IN_855 => FROM_STATE_REG_855 ,
										MUX_1024_1_IN_856 => FROM_STATE_REG_856 ,
										MUX_1024_1_IN_857 => FROM_STATE_REG_857 ,
										MUX_1024_1_IN_858 => FROM_STATE_REG_858 ,
										MUX_1024_1_IN_859 => FROM_STATE_REG_859 ,
										MUX_1024_1_IN_860 => FROM_STATE_REG_860 ,
										MUX_1024_1_IN_861 => FROM_STATE_REG_861 ,
										MUX_1024_1_IN_862 => FROM_STATE_REG_862 ,
										MUX_1024_1_IN_863 => FROM_STATE_REG_863 ,
										MUX_1024_1_IN_864 => FROM_STATE_REG_864 ,
										MUX_1024_1_IN_865 => FROM_STATE_REG_865 ,
										MUX_1024_1_IN_866 => FROM_STATE_REG_866 ,
										MUX_1024_1_IN_867 => FROM_STATE_REG_867 ,
										MUX_1024_1_IN_868 => FROM_STATE_REG_868 ,
										MUX_1024_1_IN_869 => FROM_STATE_REG_869 ,
										MUX_1024_1_IN_870 => FROM_STATE_REG_870 ,
										MUX_1024_1_IN_871 => FROM_STATE_REG_871 ,
										MUX_1024_1_IN_872 => FROM_STATE_REG_872 ,
										MUX_1024_1_IN_873 => FROM_STATE_REG_873 ,
										MUX_1024_1_IN_874 => FROM_STATE_REG_874 ,
										MUX_1024_1_IN_875 => FROM_STATE_REG_875 ,
										MUX_1024_1_IN_876 => FROM_STATE_REG_876 ,
										MUX_1024_1_IN_877 => FROM_STATE_REG_877 ,
										MUX_1024_1_IN_878 => FROM_STATE_REG_878 ,
										MUX_1024_1_IN_879 => FROM_STATE_REG_879 ,
										MUX_1024_1_IN_880 => FROM_STATE_REG_880 ,
										MUX_1024_1_IN_881 => FROM_STATE_REG_881 ,
										MUX_1024_1_IN_882 => FROM_STATE_REG_882 ,
										MUX_1024_1_IN_883 => FROM_STATE_REG_883 ,
										MUX_1024_1_IN_884 => FROM_STATE_REG_884 ,
										MUX_1024_1_IN_885 => FROM_STATE_REG_885 ,
										MUX_1024_1_IN_886 => FROM_STATE_REG_886 ,
										MUX_1024_1_IN_887 => FROM_STATE_REG_887 ,
										MUX_1024_1_IN_888 => FROM_STATE_REG_888 ,
										MUX_1024_1_IN_889 => FROM_STATE_REG_889 ,
										MUX_1024_1_IN_890 => FROM_STATE_REG_890 ,
										MUX_1024_1_IN_891 => FROM_STATE_REG_891 ,
										MUX_1024_1_IN_892 => FROM_STATE_REG_892 ,
										MUX_1024_1_IN_893 => FROM_STATE_REG_893 ,
										MUX_1024_1_IN_894 => FROM_STATE_REG_894 ,
										MUX_1024_1_IN_895 => FROM_STATE_REG_895 ,
										MUX_1024_1_IN_896 => FROM_STATE_REG_896 ,
										MUX_1024_1_IN_897 => FROM_STATE_REG_897 ,
										MUX_1024_1_IN_898 => FROM_STATE_REG_898 ,
										MUX_1024_1_IN_899 => FROM_STATE_REG_899 ,
										MUX_1024_1_IN_900 => FROM_STATE_REG_900 ,
										MUX_1024_1_IN_901 => FROM_STATE_REG_901 ,
										MUX_1024_1_IN_902 => FROM_STATE_REG_902 ,
										MUX_1024_1_IN_903 => FROM_STATE_REG_903 ,
										MUX_1024_1_IN_904 => FROM_STATE_REG_904 ,
										MUX_1024_1_IN_905 => FROM_STATE_REG_905 ,
										MUX_1024_1_IN_906 => FROM_STATE_REG_906 ,
										MUX_1024_1_IN_907 => FROM_STATE_REG_907 ,
										MUX_1024_1_IN_908 => FROM_STATE_REG_908 ,
										MUX_1024_1_IN_909 => FROM_STATE_REG_909 ,
										MUX_1024_1_IN_910 => FROM_STATE_REG_910 ,
										MUX_1024_1_IN_911 => FROM_STATE_REG_911 ,
										MUX_1024_1_IN_912 => FROM_STATE_REG_912 ,
										MUX_1024_1_IN_913 => FROM_STATE_REG_913 ,
										MUX_1024_1_IN_914 => FROM_STATE_REG_914 ,
										MUX_1024_1_IN_915 => FROM_STATE_REG_915 ,
										MUX_1024_1_IN_916 => FROM_STATE_REG_916 ,
										MUX_1024_1_IN_917 => FROM_STATE_REG_917 ,
										MUX_1024_1_IN_918 => FROM_STATE_REG_918 ,
										MUX_1024_1_IN_919 => FROM_STATE_REG_919 ,
										MUX_1024_1_IN_920 => FROM_STATE_REG_920 ,
										MUX_1024_1_IN_921 => FROM_STATE_REG_921 ,
										MUX_1024_1_IN_922 => FROM_STATE_REG_922 ,
										MUX_1024_1_IN_923 => FROM_STATE_REG_923 ,
										MUX_1024_1_IN_924 => FROM_STATE_REG_924 ,
										MUX_1024_1_IN_925 => FROM_STATE_REG_925 ,
										MUX_1024_1_IN_926 => FROM_STATE_REG_926 ,
										MUX_1024_1_IN_927 => FROM_STATE_REG_927 ,
										MUX_1024_1_IN_928 => FROM_STATE_REG_928 ,
										MUX_1024_1_IN_929 => FROM_STATE_REG_929 ,
										MUX_1024_1_IN_930 => FROM_STATE_REG_930 ,
										MUX_1024_1_IN_931 => FROM_STATE_REG_931 ,
										MUX_1024_1_IN_932 => FROM_STATE_REG_932 ,
										MUX_1024_1_IN_933 => FROM_STATE_REG_933 ,
										MUX_1024_1_IN_934 => FROM_STATE_REG_934 ,
										MUX_1024_1_IN_935 => FROM_STATE_REG_935 ,
										MUX_1024_1_IN_936 => FROM_STATE_REG_936 ,
										MUX_1024_1_IN_937 => FROM_STATE_REG_937 ,
										MUX_1024_1_IN_938 => FROM_STATE_REG_938 ,
										MUX_1024_1_IN_939 => FROM_STATE_REG_939 ,
										MUX_1024_1_IN_940 => FROM_STATE_REG_940 ,
										MUX_1024_1_IN_941 => FROM_STATE_REG_941 ,
										MUX_1024_1_IN_942 => FROM_STATE_REG_942 ,
										MUX_1024_1_IN_943 => FROM_STATE_REG_943 ,
										MUX_1024_1_IN_944 => FROM_STATE_REG_944 ,
										MUX_1024_1_IN_945 => FROM_STATE_REG_945 ,
										MUX_1024_1_IN_946 => FROM_STATE_REG_946 ,
										MUX_1024_1_IN_947 => FROM_STATE_REG_947 ,
										MUX_1024_1_IN_948 => FROM_STATE_REG_948 ,
										MUX_1024_1_IN_949 => FROM_STATE_REG_949 ,
										MUX_1024_1_IN_950 => FROM_STATE_REG_950 ,
										MUX_1024_1_IN_951 => FROM_STATE_REG_951 ,
										MUX_1024_1_IN_952 => FROM_STATE_REG_952 ,
										MUX_1024_1_IN_953 => FROM_STATE_REG_953 ,
										MUX_1024_1_IN_954 => FROM_STATE_REG_954 ,
										MUX_1024_1_IN_955 => FROM_STATE_REG_955 ,
										MUX_1024_1_IN_956 => FROM_STATE_REG_956 ,
										MUX_1024_1_IN_957 => FROM_STATE_REG_957 ,
										MUX_1024_1_IN_958 => FROM_STATE_REG_958 ,
										MUX_1024_1_IN_959 => FROM_STATE_REG_959 ,
										MUX_1024_1_IN_960 => FROM_STATE_REG_960 ,
										MUX_1024_1_IN_961 => FROM_STATE_REG_961 ,
										MUX_1024_1_IN_962 => FROM_STATE_REG_962 ,
										MUX_1024_1_IN_963 => FROM_STATE_REG_963 ,
										MUX_1024_1_IN_964 => FROM_STATE_REG_964 ,
										MUX_1024_1_IN_965 => FROM_STATE_REG_965 ,
										MUX_1024_1_IN_966 => FROM_STATE_REG_966 ,
										MUX_1024_1_IN_967 => FROM_STATE_REG_967 ,
										MUX_1024_1_IN_968 => FROM_STATE_REG_968 ,
										MUX_1024_1_IN_969 => FROM_STATE_REG_969 ,
										MUX_1024_1_IN_970 => FROM_STATE_REG_970 ,
										MUX_1024_1_IN_971 => FROM_STATE_REG_971 ,
										MUX_1024_1_IN_972 => FROM_STATE_REG_972 ,
										MUX_1024_1_IN_973 => FROM_STATE_REG_973 ,
										MUX_1024_1_IN_974 => FROM_STATE_REG_974 ,
										MUX_1024_1_IN_975 => FROM_STATE_REG_975 ,
										MUX_1024_1_IN_976 => FROM_STATE_REG_976 ,
										MUX_1024_1_IN_977 => FROM_STATE_REG_977 ,
										MUX_1024_1_IN_978 => FROM_STATE_REG_978 ,
										MUX_1024_1_IN_979 => FROM_STATE_REG_979 ,
										MUX_1024_1_IN_980 => FROM_STATE_REG_980 ,
										MUX_1024_1_IN_981 => FROM_STATE_REG_981 ,
										MUX_1024_1_IN_982 => FROM_STATE_REG_982 ,
										MUX_1024_1_IN_983 => FROM_STATE_REG_983 ,
										MUX_1024_1_IN_984 => FROM_STATE_REG_984 ,
										MUX_1024_1_IN_985 => FROM_STATE_REG_985 ,
										MUX_1024_1_IN_986 => FROM_STATE_REG_986 ,
										MUX_1024_1_IN_987 => FROM_STATE_REG_987 ,
										MUX_1024_1_IN_988 => FROM_STATE_REG_988 ,
										MUX_1024_1_IN_989 => FROM_STATE_REG_989 ,
										MUX_1024_1_IN_990 => FROM_STATE_REG_990 ,
										MUX_1024_1_IN_991 => FROM_STATE_REG_991 ,
										MUX_1024_1_IN_992 => FROM_STATE_REG_992 ,
										MUX_1024_1_IN_993 => FROM_STATE_REG_993 ,
										MUX_1024_1_IN_994 => FROM_STATE_REG_994 ,
										MUX_1024_1_IN_995 => FROM_STATE_REG_995 ,
										MUX_1024_1_IN_996 => FROM_STATE_REG_996 ,
										MUX_1024_1_IN_997 => FROM_STATE_REG_997 ,
										MUX_1024_1_IN_998 => FROM_STATE_REG_998 ,
										MUX_1024_1_IN_999 => FROM_STATE_REG_999 ,
										MUX_1024_1_IN_1000 => FROM_STATE_REG_1000 ,
										MUX_1024_1_IN_1001 => FROM_STATE_REG_1001 ,
										MUX_1024_1_IN_1002 => FROM_STATE_REG_1002 ,
										MUX_1024_1_IN_1003 => FROM_STATE_REG_1003 ,
										MUX_1024_1_IN_1004 => FROM_STATE_REG_1004 ,
										MUX_1024_1_IN_1005 => FROM_STATE_REG_1005 ,
										MUX_1024_1_IN_1006 => FROM_STATE_REG_1006 ,
										MUX_1024_1_IN_1007 => FROM_STATE_REG_1007 ,
										MUX_1024_1_IN_1008 => FROM_STATE_REG_1008 ,
										MUX_1024_1_IN_1009 => FROM_STATE_REG_1009 ,
										MUX_1024_1_IN_1010 => FROM_STATE_REG_1010 ,
										MUX_1024_1_IN_1011 => FROM_STATE_REG_1011 ,
										MUX_1024_1_IN_1012 => FROM_STATE_REG_1012 ,
										MUX_1024_1_IN_1013 => FROM_STATE_REG_1013 ,
										MUX_1024_1_IN_1014 => FROM_STATE_REG_1014 ,
										MUX_1024_1_IN_1015 => FROM_STATE_REG_1015 ,
										MUX_1024_1_IN_1016 => FROM_STATE_REG_1016 ,
										MUX_1024_1_IN_1017 => FROM_STATE_REG_1017 ,
										MUX_1024_1_IN_1018 => FROM_STATE_REG_1018 ,
										MUX_1024_1_IN_1019 => FROM_STATE_REG_1019 ,
										MUX_1024_1_IN_1020 => FROM_STATE_REG_1020 ,
										MUX_1024_1_IN_1021 => FROM_STATE_REG_1021 ,
										MUX_1024_1_IN_1022 => FROM_STATE_REG_1022 ,
										MUX_1024_1_IN_1023 => FROM_STATE_REG_1023 ,
				                    			MUX_1024_1_IN_SEL => QEP_N_10_W_0_S_0_IN_OUT_STATE_SEL ,
										MUX_1024_1_OUT_RES => SELECTED_OUTPUT
									);
MUX_REAL_IMAG_SELECTION : multiplexer_2_1 GENERIC MAP (K => K)
									PORT MAP (
										MUX_2_1_IN_0 => SELECTED_OUTPUT((2*K-1) DOWNTO K),
										MUX_2_1_IN_1 => SELECTED_OUTPUT((K-1) DOWNTO 0),
				                    			MUX_2_1_IN_SEL => QEP_N_10_W_0_S_0_IN_REAL_IMAG_SEL ,
										MUX_2_1_OUT_RES => QEP_N_10_W_0_S_0_OUT_DATA
									);

END generated;