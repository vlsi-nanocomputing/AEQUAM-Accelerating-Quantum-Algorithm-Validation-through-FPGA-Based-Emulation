LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;


ENTITY tb_control_unit IS

END ENTITY;

ARCHITECTURE behavioral OF tb_control_unit IS

	COMPONENT control_unit IS
		PORT (
			--Input signals
			CONTROL_UNIT_IN_START : IN STD_LOGIC;
			CONTROL_UNIT_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);

			--Sequential
			CONTROL_UNIT_IN_CLK : IN STD_LOGIC;
			CONTROL_UNIT_IN_CLEAR : IN STD_LOGIC;
			
			--Output signals to datapath
			CONTROL_UNIT_OUT_PIPE: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			CONTROL_UNIT_OUT_LD : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			CONTROL_UNIT_OUT_MUX_CTRL : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
			CONTROL_UNIT_OUT_SUB : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
			CONTROL_UNIT_OUT_SAVED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);

			--Done signal to enable state coefficients update
			CONTROL_UNIT_OUT_DONE : OUT STD_LOGIC);	
	END COMPONENT;

SIGNAL START, DONE, CLOCK, CLEAR : STD_LOGIC := '0';


SIGNAL OPCODE : STD_LOGIC_VECTOR (3 DOWNTO 0);

SIGNAL PIPE, LD, SAVED : STD_LOGIC_VECTOR (2 DOWNTO 0);

SIGNAL SUB : STD_LOGIC_VECTOR (1 DOWNTO 0);

SIGNAL MUX_CTRL : STD_LOGIC_VECTOR (24 DOWNTO 0);

FILE RESULT_FILE : TEXT;


BEGIN

	CLEAR <= '1', '0' AFTER 40 NS;

	CLK_GEN : PROCESS
	BEGIN
	
		--IF END_SIM = '0' THEN
		
			CLOCK <= '1';
			WAIT FOR 10 NS;
			CLOCK <= '0';
			WAIT FOR 10 NS;
		
		--ELSE
		
		--END IF;
	
	END PROCESS CLK_GEN;

	OPCODE_GEN : PROCESS(CLOCK)
		
		VARIABLE CNT : INTEGER RANGE 0 TO 12 := 0;
		--VARIABLE FINISH : STD_LOGIC := '0';
		
	BEGIN

		--START <= '0';

		IF RISING_EDGE(CLOCK) AND CLEAR = '0' THEN--AND FINISH = '0' THEN

			
			--IF CNT = 0 THEN
			
			--	START <= '1';
				--OPCODE <= (OTHERS => '0');
			
			--ELSE
				IF DONE = '1' THEN

					
					CNT := CNT + 1;
					
					IF CNT = 12 THEN
					
						--FINISH := '1';
						START <= '0';
						CNT := 0;
						
					ELSE
						START <= '1';
						
					END IF;
				ELSE 
					START <= '0';				

				END IF;
			--END IF;
			
			OPCODE <= STD_LOGIC_VECTOR(TO_UNSIGNED(CNT,4));
				
			--END_SIM <= FINISH;	
			
		ELSE
		
		END IF;


	END PROCESS OPCODE_GEN;

	DUT: control_unit 	PORT MAP (
									CONTROL_UNIT_IN_START => START ,
									CONTROL_UNIT_IN_OPCODE => OPCODE ,
									CONTROL_UNIT_IN_CLK => CLOCK ,
									CONTROL_UNIT_IN_CLEAR => CLEAR ,
									CONTROL_UNIT_OUT_PIPE => PIPE ,
									CONTROL_UNIT_OUT_LD => LD ,
									CONTROL_UNIT_OUT_MUX_CTRL => MUX_CTRL ,
									CONTROL_UNIT_OUT_SUB => SUB ,
									CONTROL_UNIT_OUT_SAVED => SAVED ,
									CONTROL_UNIT_OUT_DONE => DONE
									);

FILE_OPEN(RESULT_FILE, "ctrl_unit_res.txt", WRITE_MODE);

	SAVE_RESULTS: PROCESS(CLOCK)
	
	VARIABLE RES_LINE : LINE;
	
	BEGIN
	
		IF RISING_EDGE(CLOCK) AND CLEAR = '0' THEN
		
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(OPCODE)));

			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, PIPE);
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, LD);
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(24 DOWNTO 22))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(21 DOWNTO 20))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(19 DOWNTO 18))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(17 DOWNTO 16))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(15 DOWNTO 13))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(12 DOWNTO 11))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(10 DOWNTO 9))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(8 DOWNTO 7))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, MUX_CTRL(6));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(5 DOWNTO 3))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, TO_INTEGER(UNSIGNED(MUX_CTRL(2 DOWNTO 0))));
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, SUB);
			
			WRITE(RES_LINE, ' ');
			
			WRITE(RES_LINE, SAVED);
			
			
			WRITELINE(RESULT_FILE, RES_LINE);
		
		END IF;

	END PROCESS SAVE_RESULTS;

END behavioral;