library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_128_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_128_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_32 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_33 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_34 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_35 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_36 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_37 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_38 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_39 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_40 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_41 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_42 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_43 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_44 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_45 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_46 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_47 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_48 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_49 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_50 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_51 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_52 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_53 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_54 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_55 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_56 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_57 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_58 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_59 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_60 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_61 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_62 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_63 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_64 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_65 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_66 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_67 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_68 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_69 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_70 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_71 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_72 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_73 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_74 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_75 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_76 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_77 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_78 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_79 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_80 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_81 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_82 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_83 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_84 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_85 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_86 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_87 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_88 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_89 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_90 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_91 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_92 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_93 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_94 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_95 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_96 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_97 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_98 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_99 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_100 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_101 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_102 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_103 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_104 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_105 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_106 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_107 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_108 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_109 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_110 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_111 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_112 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_113 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_114 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_115 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_116 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_117 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_118 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_119 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_120 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_121 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_122 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_123 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_124 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_125 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_126 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_127 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_SEL : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		MUX_128_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_128_1 IS

BEGIN

	MUX_128_1_OUT_RES <= 
				MUX_128_1_IN_0 WHEN MUX_128_1_IN_SEL = "0000000" ELSE
				MUX_128_1_IN_1 WHEN MUX_128_1_IN_SEL = "0000001" ELSE
				MUX_128_1_IN_2 WHEN MUX_128_1_IN_SEL = "0000010" ELSE
				MUX_128_1_IN_3 WHEN MUX_128_1_IN_SEL = "0000011" ELSE
				MUX_128_1_IN_4 WHEN MUX_128_1_IN_SEL = "0000100" ELSE
				MUX_128_1_IN_5 WHEN MUX_128_1_IN_SEL = "0000101" ELSE
				MUX_128_1_IN_6 WHEN MUX_128_1_IN_SEL = "0000110" ELSE
				MUX_128_1_IN_7 WHEN MUX_128_1_IN_SEL = "0000111" ELSE
				MUX_128_1_IN_8 WHEN MUX_128_1_IN_SEL = "0001000" ELSE
				MUX_128_1_IN_9 WHEN MUX_128_1_IN_SEL = "0001001" ELSE
				MUX_128_1_IN_10 WHEN MUX_128_1_IN_SEL = "0001010" ELSE
				MUX_128_1_IN_11 WHEN MUX_128_1_IN_SEL = "0001011" ELSE
				MUX_128_1_IN_12 WHEN MUX_128_1_IN_SEL = "0001100" ELSE
				MUX_128_1_IN_13 WHEN MUX_128_1_IN_SEL = "0001101" ELSE
				MUX_128_1_IN_14 WHEN MUX_128_1_IN_SEL = "0001110" ELSE
				MUX_128_1_IN_15 WHEN MUX_128_1_IN_SEL = "0001111" ELSE
				MUX_128_1_IN_16 WHEN MUX_128_1_IN_SEL = "0010000" ELSE
				MUX_128_1_IN_17 WHEN MUX_128_1_IN_SEL = "0010001" ELSE
				MUX_128_1_IN_18 WHEN MUX_128_1_IN_SEL = "0010010" ELSE
				MUX_128_1_IN_19 WHEN MUX_128_1_IN_SEL = "0010011" ELSE
				MUX_128_1_IN_20 WHEN MUX_128_1_IN_SEL = "0010100" ELSE
				MUX_128_1_IN_21 WHEN MUX_128_1_IN_SEL = "0010101" ELSE
				MUX_128_1_IN_22 WHEN MUX_128_1_IN_SEL = "0010110" ELSE
				MUX_128_1_IN_23 WHEN MUX_128_1_IN_SEL = "0010111" ELSE
				MUX_128_1_IN_24 WHEN MUX_128_1_IN_SEL = "0011000" ELSE
				MUX_128_1_IN_25 WHEN MUX_128_1_IN_SEL = "0011001" ELSE
				MUX_128_1_IN_26 WHEN MUX_128_1_IN_SEL = "0011010" ELSE
				MUX_128_1_IN_27 WHEN MUX_128_1_IN_SEL = "0011011" ELSE
				MUX_128_1_IN_28 WHEN MUX_128_1_IN_SEL = "0011100" ELSE
				MUX_128_1_IN_29 WHEN MUX_128_1_IN_SEL = "0011101" ELSE
				MUX_128_1_IN_30 WHEN MUX_128_1_IN_SEL = "0011110" ELSE
				MUX_128_1_IN_31 WHEN MUX_128_1_IN_SEL = "0011111" ELSE
				MUX_128_1_IN_32 WHEN MUX_128_1_IN_SEL = "0100000" ELSE
				MUX_128_1_IN_33 WHEN MUX_128_1_IN_SEL = "0100001" ELSE
				MUX_128_1_IN_34 WHEN MUX_128_1_IN_SEL = "0100010" ELSE
				MUX_128_1_IN_35 WHEN MUX_128_1_IN_SEL = "0100011" ELSE
				MUX_128_1_IN_36 WHEN MUX_128_1_IN_SEL = "0100100" ELSE
				MUX_128_1_IN_37 WHEN MUX_128_1_IN_SEL = "0100101" ELSE
				MUX_128_1_IN_38 WHEN MUX_128_1_IN_SEL = "0100110" ELSE
				MUX_128_1_IN_39 WHEN MUX_128_1_IN_SEL = "0100111" ELSE
				MUX_128_1_IN_40 WHEN MUX_128_1_IN_SEL = "0101000" ELSE
				MUX_128_1_IN_41 WHEN MUX_128_1_IN_SEL = "0101001" ELSE
				MUX_128_1_IN_42 WHEN MUX_128_1_IN_SEL = "0101010" ELSE
				MUX_128_1_IN_43 WHEN MUX_128_1_IN_SEL = "0101011" ELSE
				MUX_128_1_IN_44 WHEN MUX_128_1_IN_SEL = "0101100" ELSE
				MUX_128_1_IN_45 WHEN MUX_128_1_IN_SEL = "0101101" ELSE
				MUX_128_1_IN_46 WHEN MUX_128_1_IN_SEL = "0101110" ELSE
				MUX_128_1_IN_47 WHEN MUX_128_1_IN_SEL = "0101111" ELSE
				MUX_128_1_IN_48 WHEN MUX_128_1_IN_SEL = "0110000" ELSE
				MUX_128_1_IN_49 WHEN MUX_128_1_IN_SEL = "0110001" ELSE
				MUX_128_1_IN_50 WHEN MUX_128_1_IN_SEL = "0110010" ELSE
				MUX_128_1_IN_51 WHEN MUX_128_1_IN_SEL = "0110011" ELSE
				MUX_128_1_IN_52 WHEN MUX_128_1_IN_SEL = "0110100" ELSE
				MUX_128_1_IN_53 WHEN MUX_128_1_IN_SEL = "0110101" ELSE
				MUX_128_1_IN_54 WHEN MUX_128_1_IN_SEL = "0110110" ELSE
				MUX_128_1_IN_55 WHEN MUX_128_1_IN_SEL = "0110111" ELSE
				MUX_128_1_IN_56 WHEN MUX_128_1_IN_SEL = "0111000" ELSE
				MUX_128_1_IN_57 WHEN MUX_128_1_IN_SEL = "0111001" ELSE
				MUX_128_1_IN_58 WHEN MUX_128_1_IN_SEL = "0111010" ELSE
				MUX_128_1_IN_59 WHEN MUX_128_1_IN_SEL = "0111011" ELSE
				MUX_128_1_IN_60 WHEN MUX_128_1_IN_SEL = "0111100" ELSE
				MUX_128_1_IN_61 WHEN MUX_128_1_IN_SEL = "0111101" ELSE
				MUX_128_1_IN_62 WHEN MUX_128_1_IN_SEL = "0111110" ELSE
				MUX_128_1_IN_63 WHEN MUX_128_1_IN_SEL = "0111111" ELSE
				MUX_128_1_IN_64 WHEN MUX_128_1_IN_SEL = "1000000" ELSE
				MUX_128_1_IN_65 WHEN MUX_128_1_IN_SEL = "1000001" ELSE
				MUX_128_1_IN_66 WHEN MUX_128_1_IN_SEL = "1000010" ELSE
				MUX_128_1_IN_67 WHEN MUX_128_1_IN_SEL = "1000011" ELSE
				MUX_128_1_IN_68 WHEN MUX_128_1_IN_SEL = "1000100" ELSE
				MUX_128_1_IN_69 WHEN MUX_128_1_IN_SEL = "1000101" ELSE
				MUX_128_1_IN_70 WHEN MUX_128_1_IN_SEL = "1000110" ELSE
				MUX_128_1_IN_71 WHEN MUX_128_1_IN_SEL = "1000111" ELSE
				MUX_128_1_IN_72 WHEN MUX_128_1_IN_SEL = "1001000" ELSE
				MUX_128_1_IN_73 WHEN MUX_128_1_IN_SEL = "1001001" ELSE
				MUX_128_1_IN_74 WHEN MUX_128_1_IN_SEL = "1001010" ELSE
				MUX_128_1_IN_75 WHEN MUX_128_1_IN_SEL = "1001011" ELSE
				MUX_128_1_IN_76 WHEN MUX_128_1_IN_SEL = "1001100" ELSE
				MUX_128_1_IN_77 WHEN MUX_128_1_IN_SEL = "1001101" ELSE
				MUX_128_1_IN_78 WHEN MUX_128_1_IN_SEL = "1001110" ELSE
				MUX_128_1_IN_79 WHEN MUX_128_1_IN_SEL = "1001111" ELSE
				MUX_128_1_IN_80 WHEN MUX_128_1_IN_SEL = "1010000" ELSE
				MUX_128_1_IN_81 WHEN MUX_128_1_IN_SEL = "1010001" ELSE
				MUX_128_1_IN_82 WHEN MUX_128_1_IN_SEL = "1010010" ELSE
				MUX_128_1_IN_83 WHEN MUX_128_1_IN_SEL = "1010011" ELSE
				MUX_128_1_IN_84 WHEN MUX_128_1_IN_SEL = "1010100" ELSE
				MUX_128_1_IN_85 WHEN MUX_128_1_IN_SEL = "1010101" ELSE
				MUX_128_1_IN_86 WHEN MUX_128_1_IN_SEL = "1010110" ELSE
				MUX_128_1_IN_87 WHEN MUX_128_1_IN_SEL = "1010111" ELSE
				MUX_128_1_IN_88 WHEN MUX_128_1_IN_SEL = "1011000" ELSE
				MUX_128_1_IN_89 WHEN MUX_128_1_IN_SEL = "1011001" ELSE
				MUX_128_1_IN_90 WHEN MUX_128_1_IN_SEL = "1011010" ELSE
				MUX_128_1_IN_91 WHEN MUX_128_1_IN_SEL = "1011011" ELSE
				MUX_128_1_IN_92 WHEN MUX_128_1_IN_SEL = "1011100" ELSE
				MUX_128_1_IN_93 WHEN MUX_128_1_IN_SEL = "1011101" ELSE
				MUX_128_1_IN_94 WHEN MUX_128_1_IN_SEL = "1011110" ELSE
				MUX_128_1_IN_95 WHEN MUX_128_1_IN_SEL = "1011111" ELSE
				MUX_128_1_IN_96 WHEN MUX_128_1_IN_SEL = "1100000" ELSE
				MUX_128_1_IN_97 WHEN MUX_128_1_IN_SEL = "1100001" ELSE
				MUX_128_1_IN_98 WHEN MUX_128_1_IN_SEL = "1100010" ELSE
				MUX_128_1_IN_99 WHEN MUX_128_1_IN_SEL = "1100011" ELSE
				MUX_128_1_IN_100 WHEN MUX_128_1_IN_SEL = "1100100" ELSE
				MUX_128_1_IN_101 WHEN MUX_128_1_IN_SEL = "1100101" ELSE
				MUX_128_1_IN_102 WHEN MUX_128_1_IN_SEL = "1100110" ELSE
				MUX_128_1_IN_103 WHEN MUX_128_1_IN_SEL = "1100111" ELSE
				MUX_128_1_IN_104 WHEN MUX_128_1_IN_SEL = "1101000" ELSE
				MUX_128_1_IN_105 WHEN MUX_128_1_IN_SEL = "1101001" ELSE
				MUX_128_1_IN_106 WHEN MUX_128_1_IN_SEL = "1101010" ELSE
				MUX_128_1_IN_107 WHEN MUX_128_1_IN_SEL = "1101011" ELSE
				MUX_128_1_IN_108 WHEN MUX_128_1_IN_SEL = "1101100" ELSE
				MUX_128_1_IN_109 WHEN MUX_128_1_IN_SEL = "1101101" ELSE
				MUX_128_1_IN_110 WHEN MUX_128_1_IN_SEL = "1101110" ELSE
				MUX_128_1_IN_111 WHEN MUX_128_1_IN_SEL = "1101111" ELSE
				MUX_128_1_IN_112 WHEN MUX_128_1_IN_SEL = "1110000" ELSE
				MUX_128_1_IN_113 WHEN MUX_128_1_IN_SEL = "1110001" ELSE
				MUX_128_1_IN_114 WHEN MUX_128_1_IN_SEL = "1110010" ELSE
				MUX_128_1_IN_115 WHEN MUX_128_1_IN_SEL = "1110011" ELSE
				MUX_128_1_IN_116 WHEN MUX_128_1_IN_SEL = "1110100" ELSE
				MUX_128_1_IN_117 WHEN MUX_128_1_IN_SEL = "1110101" ELSE
				MUX_128_1_IN_118 WHEN MUX_128_1_IN_SEL = "1110110" ELSE
				MUX_128_1_IN_119 WHEN MUX_128_1_IN_SEL = "1110111" ELSE
				MUX_128_1_IN_120 WHEN MUX_128_1_IN_SEL = "1111000" ELSE
				MUX_128_1_IN_121 WHEN MUX_128_1_IN_SEL = "1111001" ELSE
				MUX_128_1_IN_122 WHEN MUX_128_1_IN_SEL = "1111010" ELSE
				MUX_128_1_IN_123 WHEN MUX_128_1_IN_SEL = "1111011" ELSE
				MUX_128_1_IN_124 WHEN MUX_128_1_IN_SEL = "1111100" ELSE
				MUX_128_1_IN_125 WHEN MUX_128_1_IN_SEL = "1111101" ELSE
				MUX_128_1_IN_126 WHEN MUX_128_1_IN_SEL = "1111110" ELSE
				MUX_128_1_IN_127 WHEN MUX_128_1_IN_SEL = "1111111" ELSE
				(OTHERS => '0');


END behavioral;