library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_6_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_6_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		MUX_6_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_6_1 IS

BEGIN

	MUX_6_1_OUT_RES <= 
				MUX_6_1_IN_0 WHEN MUX_6_1_IN_SEL = "000" ELSE
				MUX_6_1_IN_1 WHEN MUX_6_1_IN_SEL = "001" ELSE
				MUX_6_1_IN_2 WHEN MUX_6_1_IN_SEL = "010" ELSE
				MUX_6_1_IN_3 WHEN MUX_6_1_IN_SEL = "011" ELSE
				MUX_6_1_IN_4 WHEN MUX_6_1_IN_SEL = "100" ELSE
				MUX_6_1_IN_5 WHEN MUX_6_1_IN_SEL = "101" ELSE
				(OTHERS => '0');


END behavioral;