library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_256_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_256_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_32 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_33 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_34 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_35 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_36 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_37 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_38 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_39 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_40 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_41 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_42 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_43 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_44 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_45 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_46 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_47 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_48 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_49 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_50 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_51 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_52 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_53 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_54 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_55 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_56 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_57 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_58 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_59 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_60 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_61 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_62 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_63 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_64 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_65 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_66 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_67 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_68 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_69 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_70 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_71 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_72 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_73 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_74 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_75 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_76 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_77 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_78 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_79 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_80 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_81 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_82 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_83 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_84 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_85 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_86 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_87 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_88 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_89 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_90 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_91 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_92 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_93 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_94 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_95 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_96 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_97 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_98 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_99 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_100 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_101 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_102 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_103 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_104 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_105 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_106 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_107 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_108 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_109 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_110 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_111 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_112 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_113 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_114 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_115 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_116 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_117 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_118 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_119 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_120 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_121 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_122 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_123 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_124 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_125 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_126 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_127 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_128 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_129 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_130 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_131 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_132 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_133 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_134 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_135 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_136 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_137 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_138 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_139 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_140 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_141 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_142 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_143 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_144 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_145 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_146 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_147 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_148 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_149 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_150 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_151 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_152 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_153 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_154 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_155 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_156 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_157 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_158 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_159 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_160 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_161 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_162 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_163 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_164 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_165 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_166 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_167 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_168 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_169 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_170 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_171 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_172 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_173 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_174 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_175 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_176 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_177 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_178 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_179 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_180 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_181 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_182 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_183 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_184 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_185 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_186 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_187 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_188 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_189 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_190 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_191 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_192 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_193 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_194 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_195 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_196 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_197 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_198 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_199 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_200 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_201 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_202 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_203 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_204 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_205 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_206 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_207 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_208 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_209 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_210 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_211 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_212 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_213 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_214 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_215 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_216 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_217 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_218 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_219 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_220 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_221 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_222 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_223 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_224 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_225 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_226 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_227 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_228 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_229 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_230 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_231 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_232 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_233 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_234 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_235 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_236 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_237 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_238 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_239 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_240 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_241 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_242 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_243 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_244 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_245 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_246 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_247 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_248 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_249 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_250 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_251 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_252 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_253 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_254 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_255 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_256_1_IN_SEL : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		MUX_256_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_256_1 IS

BEGIN

	MUX_256_1_OUT_RES <= 
				MUX_256_1_IN_0 WHEN MUX_256_1_IN_SEL = "00000000" ELSE
				MUX_256_1_IN_1 WHEN MUX_256_1_IN_SEL = "00000001" ELSE
				MUX_256_1_IN_2 WHEN MUX_256_1_IN_SEL = "00000010" ELSE
				MUX_256_1_IN_3 WHEN MUX_256_1_IN_SEL = "00000011" ELSE
				MUX_256_1_IN_4 WHEN MUX_256_1_IN_SEL = "00000100" ELSE
				MUX_256_1_IN_5 WHEN MUX_256_1_IN_SEL = "00000101" ELSE
				MUX_256_1_IN_6 WHEN MUX_256_1_IN_SEL = "00000110" ELSE
				MUX_256_1_IN_7 WHEN MUX_256_1_IN_SEL = "00000111" ELSE
				MUX_256_1_IN_8 WHEN MUX_256_1_IN_SEL = "00001000" ELSE
				MUX_256_1_IN_9 WHEN MUX_256_1_IN_SEL = "00001001" ELSE
				MUX_256_1_IN_10 WHEN MUX_256_1_IN_SEL = "00001010" ELSE
				MUX_256_1_IN_11 WHEN MUX_256_1_IN_SEL = "00001011" ELSE
				MUX_256_1_IN_12 WHEN MUX_256_1_IN_SEL = "00001100" ELSE
				MUX_256_1_IN_13 WHEN MUX_256_1_IN_SEL = "00001101" ELSE
				MUX_256_1_IN_14 WHEN MUX_256_1_IN_SEL = "00001110" ELSE
				MUX_256_1_IN_15 WHEN MUX_256_1_IN_SEL = "00001111" ELSE
				MUX_256_1_IN_16 WHEN MUX_256_1_IN_SEL = "00010000" ELSE
				MUX_256_1_IN_17 WHEN MUX_256_1_IN_SEL = "00010001" ELSE
				MUX_256_1_IN_18 WHEN MUX_256_1_IN_SEL = "00010010" ELSE
				MUX_256_1_IN_19 WHEN MUX_256_1_IN_SEL = "00010011" ELSE
				MUX_256_1_IN_20 WHEN MUX_256_1_IN_SEL = "00010100" ELSE
				MUX_256_1_IN_21 WHEN MUX_256_1_IN_SEL = "00010101" ELSE
				MUX_256_1_IN_22 WHEN MUX_256_1_IN_SEL = "00010110" ELSE
				MUX_256_1_IN_23 WHEN MUX_256_1_IN_SEL = "00010111" ELSE
				MUX_256_1_IN_24 WHEN MUX_256_1_IN_SEL = "00011000" ELSE
				MUX_256_1_IN_25 WHEN MUX_256_1_IN_SEL = "00011001" ELSE
				MUX_256_1_IN_26 WHEN MUX_256_1_IN_SEL = "00011010" ELSE
				MUX_256_1_IN_27 WHEN MUX_256_1_IN_SEL = "00011011" ELSE
				MUX_256_1_IN_28 WHEN MUX_256_1_IN_SEL = "00011100" ELSE
				MUX_256_1_IN_29 WHEN MUX_256_1_IN_SEL = "00011101" ELSE
				MUX_256_1_IN_30 WHEN MUX_256_1_IN_SEL = "00011110" ELSE
				MUX_256_1_IN_31 WHEN MUX_256_1_IN_SEL = "00011111" ELSE
				MUX_256_1_IN_32 WHEN MUX_256_1_IN_SEL = "00100000" ELSE
				MUX_256_1_IN_33 WHEN MUX_256_1_IN_SEL = "00100001" ELSE
				MUX_256_1_IN_34 WHEN MUX_256_1_IN_SEL = "00100010" ELSE
				MUX_256_1_IN_35 WHEN MUX_256_1_IN_SEL = "00100011" ELSE
				MUX_256_1_IN_36 WHEN MUX_256_1_IN_SEL = "00100100" ELSE
				MUX_256_1_IN_37 WHEN MUX_256_1_IN_SEL = "00100101" ELSE
				MUX_256_1_IN_38 WHEN MUX_256_1_IN_SEL = "00100110" ELSE
				MUX_256_1_IN_39 WHEN MUX_256_1_IN_SEL = "00100111" ELSE
				MUX_256_1_IN_40 WHEN MUX_256_1_IN_SEL = "00101000" ELSE
				MUX_256_1_IN_41 WHEN MUX_256_1_IN_SEL = "00101001" ELSE
				MUX_256_1_IN_42 WHEN MUX_256_1_IN_SEL = "00101010" ELSE
				MUX_256_1_IN_43 WHEN MUX_256_1_IN_SEL = "00101011" ELSE
				MUX_256_1_IN_44 WHEN MUX_256_1_IN_SEL = "00101100" ELSE
				MUX_256_1_IN_45 WHEN MUX_256_1_IN_SEL = "00101101" ELSE
				MUX_256_1_IN_46 WHEN MUX_256_1_IN_SEL = "00101110" ELSE
				MUX_256_1_IN_47 WHEN MUX_256_1_IN_SEL = "00101111" ELSE
				MUX_256_1_IN_48 WHEN MUX_256_1_IN_SEL = "00110000" ELSE
				MUX_256_1_IN_49 WHEN MUX_256_1_IN_SEL = "00110001" ELSE
				MUX_256_1_IN_50 WHEN MUX_256_1_IN_SEL = "00110010" ELSE
				MUX_256_1_IN_51 WHEN MUX_256_1_IN_SEL = "00110011" ELSE
				MUX_256_1_IN_52 WHEN MUX_256_1_IN_SEL = "00110100" ELSE
				MUX_256_1_IN_53 WHEN MUX_256_1_IN_SEL = "00110101" ELSE
				MUX_256_1_IN_54 WHEN MUX_256_1_IN_SEL = "00110110" ELSE
				MUX_256_1_IN_55 WHEN MUX_256_1_IN_SEL = "00110111" ELSE
				MUX_256_1_IN_56 WHEN MUX_256_1_IN_SEL = "00111000" ELSE
				MUX_256_1_IN_57 WHEN MUX_256_1_IN_SEL = "00111001" ELSE
				MUX_256_1_IN_58 WHEN MUX_256_1_IN_SEL = "00111010" ELSE
				MUX_256_1_IN_59 WHEN MUX_256_1_IN_SEL = "00111011" ELSE
				MUX_256_1_IN_60 WHEN MUX_256_1_IN_SEL = "00111100" ELSE
				MUX_256_1_IN_61 WHEN MUX_256_1_IN_SEL = "00111101" ELSE
				MUX_256_1_IN_62 WHEN MUX_256_1_IN_SEL = "00111110" ELSE
				MUX_256_1_IN_63 WHEN MUX_256_1_IN_SEL = "00111111" ELSE
				MUX_256_1_IN_64 WHEN MUX_256_1_IN_SEL = "01000000" ELSE
				MUX_256_1_IN_65 WHEN MUX_256_1_IN_SEL = "01000001" ELSE
				MUX_256_1_IN_66 WHEN MUX_256_1_IN_SEL = "01000010" ELSE
				MUX_256_1_IN_67 WHEN MUX_256_1_IN_SEL = "01000011" ELSE
				MUX_256_1_IN_68 WHEN MUX_256_1_IN_SEL = "01000100" ELSE
				MUX_256_1_IN_69 WHEN MUX_256_1_IN_SEL = "01000101" ELSE
				MUX_256_1_IN_70 WHEN MUX_256_1_IN_SEL = "01000110" ELSE
				MUX_256_1_IN_71 WHEN MUX_256_1_IN_SEL = "01000111" ELSE
				MUX_256_1_IN_72 WHEN MUX_256_1_IN_SEL = "01001000" ELSE
				MUX_256_1_IN_73 WHEN MUX_256_1_IN_SEL = "01001001" ELSE
				MUX_256_1_IN_74 WHEN MUX_256_1_IN_SEL = "01001010" ELSE
				MUX_256_1_IN_75 WHEN MUX_256_1_IN_SEL = "01001011" ELSE
				MUX_256_1_IN_76 WHEN MUX_256_1_IN_SEL = "01001100" ELSE
				MUX_256_1_IN_77 WHEN MUX_256_1_IN_SEL = "01001101" ELSE
				MUX_256_1_IN_78 WHEN MUX_256_1_IN_SEL = "01001110" ELSE
				MUX_256_1_IN_79 WHEN MUX_256_1_IN_SEL = "01001111" ELSE
				MUX_256_1_IN_80 WHEN MUX_256_1_IN_SEL = "01010000" ELSE
				MUX_256_1_IN_81 WHEN MUX_256_1_IN_SEL = "01010001" ELSE
				MUX_256_1_IN_82 WHEN MUX_256_1_IN_SEL = "01010010" ELSE
				MUX_256_1_IN_83 WHEN MUX_256_1_IN_SEL = "01010011" ELSE
				MUX_256_1_IN_84 WHEN MUX_256_1_IN_SEL = "01010100" ELSE
				MUX_256_1_IN_85 WHEN MUX_256_1_IN_SEL = "01010101" ELSE
				MUX_256_1_IN_86 WHEN MUX_256_1_IN_SEL = "01010110" ELSE
				MUX_256_1_IN_87 WHEN MUX_256_1_IN_SEL = "01010111" ELSE
				MUX_256_1_IN_88 WHEN MUX_256_1_IN_SEL = "01011000" ELSE
				MUX_256_1_IN_89 WHEN MUX_256_1_IN_SEL = "01011001" ELSE
				MUX_256_1_IN_90 WHEN MUX_256_1_IN_SEL = "01011010" ELSE
				MUX_256_1_IN_91 WHEN MUX_256_1_IN_SEL = "01011011" ELSE
				MUX_256_1_IN_92 WHEN MUX_256_1_IN_SEL = "01011100" ELSE
				MUX_256_1_IN_93 WHEN MUX_256_1_IN_SEL = "01011101" ELSE
				MUX_256_1_IN_94 WHEN MUX_256_1_IN_SEL = "01011110" ELSE
				MUX_256_1_IN_95 WHEN MUX_256_1_IN_SEL = "01011111" ELSE
				MUX_256_1_IN_96 WHEN MUX_256_1_IN_SEL = "01100000" ELSE
				MUX_256_1_IN_97 WHEN MUX_256_1_IN_SEL = "01100001" ELSE
				MUX_256_1_IN_98 WHEN MUX_256_1_IN_SEL = "01100010" ELSE
				MUX_256_1_IN_99 WHEN MUX_256_1_IN_SEL = "01100011" ELSE
				MUX_256_1_IN_100 WHEN MUX_256_1_IN_SEL = "01100100" ELSE
				MUX_256_1_IN_101 WHEN MUX_256_1_IN_SEL = "01100101" ELSE
				MUX_256_1_IN_102 WHEN MUX_256_1_IN_SEL = "01100110" ELSE
				MUX_256_1_IN_103 WHEN MUX_256_1_IN_SEL = "01100111" ELSE
				MUX_256_1_IN_104 WHEN MUX_256_1_IN_SEL = "01101000" ELSE
				MUX_256_1_IN_105 WHEN MUX_256_1_IN_SEL = "01101001" ELSE
				MUX_256_1_IN_106 WHEN MUX_256_1_IN_SEL = "01101010" ELSE
				MUX_256_1_IN_107 WHEN MUX_256_1_IN_SEL = "01101011" ELSE
				MUX_256_1_IN_108 WHEN MUX_256_1_IN_SEL = "01101100" ELSE
				MUX_256_1_IN_109 WHEN MUX_256_1_IN_SEL = "01101101" ELSE
				MUX_256_1_IN_110 WHEN MUX_256_1_IN_SEL = "01101110" ELSE
				MUX_256_1_IN_111 WHEN MUX_256_1_IN_SEL = "01101111" ELSE
				MUX_256_1_IN_112 WHEN MUX_256_1_IN_SEL = "01110000" ELSE
				MUX_256_1_IN_113 WHEN MUX_256_1_IN_SEL = "01110001" ELSE
				MUX_256_1_IN_114 WHEN MUX_256_1_IN_SEL = "01110010" ELSE
				MUX_256_1_IN_115 WHEN MUX_256_1_IN_SEL = "01110011" ELSE
				MUX_256_1_IN_116 WHEN MUX_256_1_IN_SEL = "01110100" ELSE
				MUX_256_1_IN_117 WHEN MUX_256_1_IN_SEL = "01110101" ELSE
				MUX_256_1_IN_118 WHEN MUX_256_1_IN_SEL = "01110110" ELSE
				MUX_256_1_IN_119 WHEN MUX_256_1_IN_SEL = "01110111" ELSE
				MUX_256_1_IN_120 WHEN MUX_256_1_IN_SEL = "01111000" ELSE
				MUX_256_1_IN_121 WHEN MUX_256_1_IN_SEL = "01111001" ELSE
				MUX_256_1_IN_122 WHEN MUX_256_1_IN_SEL = "01111010" ELSE
				MUX_256_1_IN_123 WHEN MUX_256_1_IN_SEL = "01111011" ELSE
				MUX_256_1_IN_124 WHEN MUX_256_1_IN_SEL = "01111100" ELSE
				MUX_256_1_IN_125 WHEN MUX_256_1_IN_SEL = "01111101" ELSE
				MUX_256_1_IN_126 WHEN MUX_256_1_IN_SEL = "01111110" ELSE
				MUX_256_1_IN_127 WHEN MUX_256_1_IN_SEL = "01111111" ELSE
				MUX_256_1_IN_128 WHEN MUX_256_1_IN_SEL = "10000000" ELSE
				MUX_256_1_IN_129 WHEN MUX_256_1_IN_SEL = "10000001" ELSE
				MUX_256_1_IN_130 WHEN MUX_256_1_IN_SEL = "10000010" ELSE
				MUX_256_1_IN_131 WHEN MUX_256_1_IN_SEL = "10000011" ELSE
				MUX_256_1_IN_132 WHEN MUX_256_1_IN_SEL = "10000100" ELSE
				MUX_256_1_IN_133 WHEN MUX_256_1_IN_SEL = "10000101" ELSE
				MUX_256_1_IN_134 WHEN MUX_256_1_IN_SEL = "10000110" ELSE
				MUX_256_1_IN_135 WHEN MUX_256_1_IN_SEL = "10000111" ELSE
				MUX_256_1_IN_136 WHEN MUX_256_1_IN_SEL = "10001000" ELSE
				MUX_256_1_IN_137 WHEN MUX_256_1_IN_SEL = "10001001" ELSE
				MUX_256_1_IN_138 WHEN MUX_256_1_IN_SEL = "10001010" ELSE
				MUX_256_1_IN_139 WHEN MUX_256_1_IN_SEL = "10001011" ELSE
				MUX_256_1_IN_140 WHEN MUX_256_1_IN_SEL = "10001100" ELSE
				MUX_256_1_IN_141 WHEN MUX_256_1_IN_SEL = "10001101" ELSE
				MUX_256_1_IN_142 WHEN MUX_256_1_IN_SEL = "10001110" ELSE
				MUX_256_1_IN_143 WHEN MUX_256_1_IN_SEL = "10001111" ELSE
				MUX_256_1_IN_144 WHEN MUX_256_1_IN_SEL = "10010000" ELSE
				MUX_256_1_IN_145 WHEN MUX_256_1_IN_SEL = "10010001" ELSE
				MUX_256_1_IN_146 WHEN MUX_256_1_IN_SEL = "10010010" ELSE
				MUX_256_1_IN_147 WHEN MUX_256_1_IN_SEL = "10010011" ELSE
				MUX_256_1_IN_148 WHEN MUX_256_1_IN_SEL = "10010100" ELSE
				MUX_256_1_IN_149 WHEN MUX_256_1_IN_SEL = "10010101" ELSE
				MUX_256_1_IN_150 WHEN MUX_256_1_IN_SEL = "10010110" ELSE
				MUX_256_1_IN_151 WHEN MUX_256_1_IN_SEL = "10010111" ELSE
				MUX_256_1_IN_152 WHEN MUX_256_1_IN_SEL = "10011000" ELSE
				MUX_256_1_IN_153 WHEN MUX_256_1_IN_SEL = "10011001" ELSE
				MUX_256_1_IN_154 WHEN MUX_256_1_IN_SEL = "10011010" ELSE
				MUX_256_1_IN_155 WHEN MUX_256_1_IN_SEL = "10011011" ELSE
				MUX_256_1_IN_156 WHEN MUX_256_1_IN_SEL = "10011100" ELSE
				MUX_256_1_IN_157 WHEN MUX_256_1_IN_SEL = "10011101" ELSE
				MUX_256_1_IN_158 WHEN MUX_256_1_IN_SEL = "10011110" ELSE
				MUX_256_1_IN_159 WHEN MUX_256_1_IN_SEL = "10011111" ELSE
				MUX_256_1_IN_160 WHEN MUX_256_1_IN_SEL = "10100000" ELSE
				MUX_256_1_IN_161 WHEN MUX_256_1_IN_SEL = "10100001" ELSE
				MUX_256_1_IN_162 WHEN MUX_256_1_IN_SEL = "10100010" ELSE
				MUX_256_1_IN_163 WHEN MUX_256_1_IN_SEL = "10100011" ELSE
				MUX_256_1_IN_164 WHEN MUX_256_1_IN_SEL = "10100100" ELSE
				MUX_256_1_IN_165 WHEN MUX_256_1_IN_SEL = "10100101" ELSE
				MUX_256_1_IN_166 WHEN MUX_256_1_IN_SEL = "10100110" ELSE
				MUX_256_1_IN_167 WHEN MUX_256_1_IN_SEL = "10100111" ELSE
				MUX_256_1_IN_168 WHEN MUX_256_1_IN_SEL = "10101000" ELSE
				MUX_256_1_IN_169 WHEN MUX_256_1_IN_SEL = "10101001" ELSE
				MUX_256_1_IN_170 WHEN MUX_256_1_IN_SEL = "10101010" ELSE
				MUX_256_1_IN_171 WHEN MUX_256_1_IN_SEL = "10101011" ELSE
				MUX_256_1_IN_172 WHEN MUX_256_1_IN_SEL = "10101100" ELSE
				MUX_256_1_IN_173 WHEN MUX_256_1_IN_SEL = "10101101" ELSE
				MUX_256_1_IN_174 WHEN MUX_256_1_IN_SEL = "10101110" ELSE
				MUX_256_1_IN_175 WHEN MUX_256_1_IN_SEL = "10101111" ELSE
				MUX_256_1_IN_176 WHEN MUX_256_1_IN_SEL = "10110000" ELSE
				MUX_256_1_IN_177 WHEN MUX_256_1_IN_SEL = "10110001" ELSE
				MUX_256_1_IN_178 WHEN MUX_256_1_IN_SEL = "10110010" ELSE
				MUX_256_1_IN_179 WHEN MUX_256_1_IN_SEL = "10110011" ELSE
				MUX_256_1_IN_180 WHEN MUX_256_1_IN_SEL = "10110100" ELSE
				MUX_256_1_IN_181 WHEN MUX_256_1_IN_SEL = "10110101" ELSE
				MUX_256_1_IN_182 WHEN MUX_256_1_IN_SEL = "10110110" ELSE
				MUX_256_1_IN_183 WHEN MUX_256_1_IN_SEL = "10110111" ELSE
				MUX_256_1_IN_184 WHEN MUX_256_1_IN_SEL = "10111000" ELSE
				MUX_256_1_IN_185 WHEN MUX_256_1_IN_SEL = "10111001" ELSE
				MUX_256_1_IN_186 WHEN MUX_256_1_IN_SEL = "10111010" ELSE
				MUX_256_1_IN_187 WHEN MUX_256_1_IN_SEL = "10111011" ELSE
				MUX_256_1_IN_188 WHEN MUX_256_1_IN_SEL = "10111100" ELSE
				MUX_256_1_IN_189 WHEN MUX_256_1_IN_SEL = "10111101" ELSE
				MUX_256_1_IN_190 WHEN MUX_256_1_IN_SEL = "10111110" ELSE
				MUX_256_1_IN_191 WHEN MUX_256_1_IN_SEL = "10111111" ELSE
				MUX_256_1_IN_192 WHEN MUX_256_1_IN_SEL = "11000000" ELSE
				MUX_256_1_IN_193 WHEN MUX_256_1_IN_SEL = "11000001" ELSE
				MUX_256_1_IN_194 WHEN MUX_256_1_IN_SEL = "11000010" ELSE
				MUX_256_1_IN_195 WHEN MUX_256_1_IN_SEL = "11000011" ELSE
				MUX_256_1_IN_196 WHEN MUX_256_1_IN_SEL = "11000100" ELSE
				MUX_256_1_IN_197 WHEN MUX_256_1_IN_SEL = "11000101" ELSE
				MUX_256_1_IN_198 WHEN MUX_256_1_IN_SEL = "11000110" ELSE
				MUX_256_1_IN_199 WHEN MUX_256_1_IN_SEL = "11000111" ELSE
				MUX_256_1_IN_200 WHEN MUX_256_1_IN_SEL = "11001000" ELSE
				MUX_256_1_IN_201 WHEN MUX_256_1_IN_SEL = "11001001" ELSE
				MUX_256_1_IN_202 WHEN MUX_256_1_IN_SEL = "11001010" ELSE
				MUX_256_1_IN_203 WHEN MUX_256_1_IN_SEL = "11001011" ELSE
				MUX_256_1_IN_204 WHEN MUX_256_1_IN_SEL = "11001100" ELSE
				MUX_256_1_IN_205 WHEN MUX_256_1_IN_SEL = "11001101" ELSE
				MUX_256_1_IN_206 WHEN MUX_256_1_IN_SEL = "11001110" ELSE
				MUX_256_1_IN_207 WHEN MUX_256_1_IN_SEL = "11001111" ELSE
				MUX_256_1_IN_208 WHEN MUX_256_1_IN_SEL = "11010000" ELSE
				MUX_256_1_IN_209 WHEN MUX_256_1_IN_SEL = "11010001" ELSE
				MUX_256_1_IN_210 WHEN MUX_256_1_IN_SEL = "11010010" ELSE
				MUX_256_1_IN_211 WHEN MUX_256_1_IN_SEL = "11010011" ELSE
				MUX_256_1_IN_212 WHEN MUX_256_1_IN_SEL = "11010100" ELSE
				MUX_256_1_IN_213 WHEN MUX_256_1_IN_SEL = "11010101" ELSE
				MUX_256_1_IN_214 WHEN MUX_256_1_IN_SEL = "11010110" ELSE
				MUX_256_1_IN_215 WHEN MUX_256_1_IN_SEL = "11010111" ELSE
				MUX_256_1_IN_216 WHEN MUX_256_1_IN_SEL = "11011000" ELSE
				MUX_256_1_IN_217 WHEN MUX_256_1_IN_SEL = "11011001" ELSE
				MUX_256_1_IN_218 WHEN MUX_256_1_IN_SEL = "11011010" ELSE
				MUX_256_1_IN_219 WHEN MUX_256_1_IN_SEL = "11011011" ELSE
				MUX_256_1_IN_220 WHEN MUX_256_1_IN_SEL = "11011100" ELSE
				MUX_256_1_IN_221 WHEN MUX_256_1_IN_SEL = "11011101" ELSE
				MUX_256_1_IN_222 WHEN MUX_256_1_IN_SEL = "11011110" ELSE
				MUX_256_1_IN_223 WHEN MUX_256_1_IN_SEL = "11011111" ELSE
				MUX_256_1_IN_224 WHEN MUX_256_1_IN_SEL = "11100000" ELSE
				MUX_256_1_IN_225 WHEN MUX_256_1_IN_SEL = "11100001" ELSE
				MUX_256_1_IN_226 WHEN MUX_256_1_IN_SEL = "11100010" ELSE
				MUX_256_1_IN_227 WHEN MUX_256_1_IN_SEL = "11100011" ELSE
				MUX_256_1_IN_228 WHEN MUX_256_1_IN_SEL = "11100100" ELSE
				MUX_256_1_IN_229 WHEN MUX_256_1_IN_SEL = "11100101" ELSE
				MUX_256_1_IN_230 WHEN MUX_256_1_IN_SEL = "11100110" ELSE
				MUX_256_1_IN_231 WHEN MUX_256_1_IN_SEL = "11100111" ELSE
				MUX_256_1_IN_232 WHEN MUX_256_1_IN_SEL = "11101000" ELSE
				MUX_256_1_IN_233 WHEN MUX_256_1_IN_SEL = "11101001" ELSE
				MUX_256_1_IN_234 WHEN MUX_256_1_IN_SEL = "11101010" ELSE
				MUX_256_1_IN_235 WHEN MUX_256_1_IN_SEL = "11101011" ELSE
				MUX_256_1_IN_236 WHEN MUX_256_1_IN_SEL = "11101100" ELSE
				MUX_256_1_IN_237 WHEN MUX_256_1_IN_SEL = "11101101" ELSE
				MUX_256_1_IN_238 WHEN MUX_256_1_IN_SEL = "11101110" ELSE
				MUX_256_1_IN_239 WHEN MUX_256_1_IN_SEL = "11101111" ELSE
				MUX_256_1_IN_240 WHEN MUX_256_1_IN_SEL = "11110000" ELSE
				MUX_256_1_IN_241 WHEN MUX_256_1_IN_SEL = "11110001" ELSE
				MUX_256_1_IN_242 WHEN MUX_256_1_IN_SEL = "11110010" ELSE
				MUX_256_1_IN_243 WHEN MUX_256_1_IN_SEL = "11110011" ELSE
				MUX_256_1_IN_244 WHEN MUX_256_1_IN_SEL = "11110100" ELSE
				MUX_256_1_IN_245 WHEN MUX_256_1_IN_SEL = "11110101" ELSE
				MUX_256_1_IN_246 WHEN MUX_256_1_IN_SEL = "11110110" ELSE
				MUX_256_1_IN_247 WHEN MUX_256_1_IN_SEL = "11110111" ELSE
				MUX_256_1_IN_248 WHEN MUX_256_1_IN_SEL = "11111000" ELSE
				MUX_256_1_IN_249 WHEN MUX_256_1_IN_SEL = "11111001" ELSE
				MUX_256_1_IN_250 WHEN MUX_256_1_IN_SEL = "11111010" ELSE
				MUX_256_1_IN_251 WHEN MUX_256_1_IN_SEL = "11111011" ELSE
				MUX_256_1_IN_252 WHEN MUX_256_1_IN_SEL = "11111100" ELSE
				MUX_256_1_IN_253 WHEN MUX_256_1_IN_SEL = "11111101" ELSE
				MUX_256_1_IN_254 WHEN MUX_256_1_IN_SEL = "11111110" ELSE
				MUX_256_1_IN_255 WHEN MUX_256_1_IN_SEL = "11111111" ELSE
				(OTHERS => '0');


END behavioral;