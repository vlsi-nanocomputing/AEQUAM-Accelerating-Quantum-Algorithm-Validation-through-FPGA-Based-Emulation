library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY QEP_N_7_W_5_S_0 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		QEP_N_7_W_5_S_0_IN_START : IN STD_LOGIC;
		QEP_N_7_W_5_S_0_IN_QTGT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);  
		QEP_N_7_W_5_S_0_IN_CTRL_MASK : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		QEP_N_7_W_5_S_0_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		QEP_N_7_W_5_S_0_IN_SIN : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_7_W_5_S_0_IN_COS : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_7_W_5_S_0_IN_WIN_SEL : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		QEP_N_7_W_5_S_0_IN_OUT_STATE_SEL : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		QEP_N_7_W_5_S_0_IN_REAL_IMAG_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		QEP_N_7_W_5_S_0_IN_CLK : IN STD_LOGIC;
		QEP_N_7_W_5_S_0_IN_CLEAR : IN STD_LOGIC;
		QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF : IN STD_LOGIC;
		QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE : IN STD_LOGIC;
		QEP_N_7_W_5_S_0_OUT_DONE : OUT STD_LOGIC;
		QEP_N_7_W_5_S_0_OUT_DATA : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;
ARCHITECTURE generated OF QEP_N_7_W_5_S_0 IS
COMPONENT multiplexer_2_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_2_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		MUX_2_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_7_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_7_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_7_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_7_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_7_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_7_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_7_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_7_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_7_1_IN_SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		MUX_7_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_128_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_128_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_32 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_33 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_34 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_35 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_36 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_37 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_38 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_39 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_40 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_41 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_42 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_43 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_44 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_45 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_46 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_47 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_48 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_49 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_50 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_51 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_52 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_53 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_54 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_55 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_56 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_57 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_58 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_59 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_60 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_61 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_62 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_63 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_64 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_65 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_66 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_67 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_68 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_69 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_70 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_71 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_72 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_73 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_74 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_75 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_76 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_77 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_78 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_79 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_80 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_81 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_82 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_83 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_84 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_85 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_86 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_87 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_88 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_89 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_90 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_91 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_92 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_93 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_94 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_95 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_96 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_97 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_98 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_99 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_100 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_101 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_102 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_103 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_104 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_105 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_106 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_107 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_108 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_109 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_110 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_111 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_112 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_113 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_114 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_115 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_116 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_117 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_118 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_119 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_120 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_121 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_122 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_123 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_124 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_125 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_126 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_127 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_128_1_IN_SEL : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		MUX_128_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_32_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_32_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_SEL : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		MUX_32_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register_clear_1 IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT datapath is
    GENERIC (K : INTEGER := 20);	--K represents the chosen parallelism
	PORT(
		--Data signals
		DATAPATH_IN_A : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_B : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_SINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_COSINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_PIPE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_LD : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_MUX_CTRL : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
		DATAPATH_IN_SUB : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		DATAPATH_IN_SAVED : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_CLEAR : IN STD_LOGIC;
		DATAPATH_IN_CLK : IN STD_LOGIC;
		DATAPATH_OUT_A : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_OUT_B : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0));
END COMPONENT;
COMPONENT control_unit IS
 	PORT (
		--Input signals
		CONTROL_UNIT_IN_START : IN STD_LOGIC;
		CONTROL_UNIT_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CONTROL_UNIT_IN_CLK : IN STD_LOGIC;
		CONTROL_UNIT_IN_CLEAR : IN STD_LOGIC;
		CONTROL_UNIT_OUT_PIPE: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_LD : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_MUX_CTRL : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
		CONTROL_UNIT_OUT_SUB : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		CONTROL_UNIT_OUT_SAVED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_DONE : OUT STD_LOGIC);
END COMPONENT;

SIGNAL TO_STATE_REG_0,TO_STATE_REG_1,TO_STATE_REG_2,TO_STATE_REG_3,TO_STATE_REG_4,TO_STATE_REG_5,TO_STATE_REG_6,TO_STATE_REG_7,TO_STATE_REG_8,TO_STATE_REG_9,TO_STATE_REG_10,TO_STATE_REG_11,TO_STATE_REG_12,TO_STATE_REG_13,TO_STATE_REG_14,TO_STATE_REG_15,TO_STATE_REG_16,TO_STATE_REG_17,TO_STATE_REG_18,TO_STATE_REG_19,TO_STATE_REG_20,TO_STATE_REG_21,TO_STATE_REG_22,TO_STATE_REG_23,TO_STATE_REG_24,TO_STATE_REG_25,TO_STATE_REG_26,TO_STATE_REG_27,TO_STATE_REG_28,TO_STATE_REG_29,TO_STATE_REG_30,TO_STATE_REG_31,TO_STATE_REG_32,TO_STATE_REG_33,TO_STATE_REG_34,TO_STATE_REG_35,TO_STATE_REG_36,TO_STATE_REG_37,TO_STATE_REG_38,TO_STATE_REG_39,TO_STATE_REG_40,TO_STATE_REG_41,TO_STATE_REG_42,TO_STATE_REG_43,TO_STATE_REG_44,TO_STATE_REG_45,TO_STATE_REG_46,TO_STATE_REG_47,TO_STATE_REG_48,TO_STATE_REG_49,TO_STATE_REG_50,TO_STATE_REG_51,TO_STATE_REG_52,TO_STATE_REG_53,TO_STATE_REG_54,TO_STATE_REG_55,TO_STATE_REG_56,TO_STATE_REG_57,TO_STATE_REG_58,TO_STATE_REG_59,TO_STATE_REG_60,TO_STATE_REG_61,TO_STATE_REG_62,TO_STATE_REG_63,TO_STATE_REG_64,TO_STATE_REG_65,TO_STATE_REG_66,TO_STATE_REG_67,TO_STATE_REG_68,TO_STATE_REG_69,TO_STATE_REG_70,TO_STATE_REG_71,TO_STATE_REG_72,TO_STATE_REG_73,TO_STATE_REG_74,TO_STATE_REG_75,TO_STATE_REG_76,TO_STATE_REG_77,TO_STATE_REG_78,TO_STATE_REG_79,TO_STATE_REG_80,TO_STATE_REG_81,TO_STATE_REG_82,TO_STATE_REG_83,TO_STATE_REG_84,TO_STATE_REG_85,TO_STATE_REG_86,TO_STATE_REG_87,TO_STATE_REG_88,TO_STATE_REG_89,TO_STATE_REG_90,TO_STATE_REG_91,TO_STATE_REG_92,TO_STATE_REG_93,TO_STATE_REG_94,TO_STATE_REG_95,TO_STATE_REG_96,TO_STATE_REG_97,TO_STATE_REG_98,TO_STATE_REG_99,TO_STATE_REG_100,TO_STATE_REG_101,TO_STATE_REG_102,TO_STATE_REG_103,TO_STATE_REG_104,TO_STATE_REG_105,TO_STATE_REG_106,TO_STATE_REG_107,TO_STATE_REG_108,TO_STATE_REG_109,TO_STATE_REG_110,TO_STATE_REG_111,TO_STATE_REG_112,TO_STATE_REG_113,TO_STATE_REG_114,TO_STATE_REG_115,TO_STATE_REG_116,TO_STATE_REG_117,TO_STATE_REG_118,TO_STATE_REG_119,TO_STATE_REG_120,TO_STATE_REG_121,TO_STATE_REG_122,TO_STATE_REG_123,TO_STATE_REG_124,TO_STATE_REG_125,TO_STATE_REG_126,TO_STATE_REG_127: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_STATE_REG_0,FROM_STATE_REG_1,FROM_STATE_REG_2,FROM_STATE_REG_3,FROM_STATE_REG_4,FROM_STATE_REG_5,FROM_STATE_REG_6,FROM_STATE_REG_7,FROM_STATE_REG_8,FROM_STATE_REG_9,FROM_STATE_REG_10,FROM_STATE_REG_11,FROM_STATE_REG_12,FROM_STATE_REG_13,FROM_STATE_REG_14,FROM_STATE_REG_15,FROM_STATE_REG_16,FROM_STATE_REG_17,FROM_STATE_REG_18,FROM_STATE_REG_19,FROM_STATE_REG_20,FROM_STATE_REG_21,FROM_STATE_REG_22,FROM_STATE_REG_23,FROM_STATE_REG_24,FROM_STATE_REG_25,FROM_STATE_REG_26,FROM_STATE_REG_27,FROM_STATE_REG_28,FROM_STATE_REG_29,FROM_STATE_REG_30,FROM_STATE_REG_31,FROM_STATE_REG_32,FROM_STATE_REG_33,FROM_STATE_REG_34,FROM_STATE_REG_35,FROM_STATE_REG_36,FROM_STATE_REG_37,FROM_STATE_REG_38,FROM_STATE_REG_39,FROM_STATE_REG_40,FROM_STATE_REG_41,FROM_STATE_REG_42,FROM_STATE_REG_43,FROM_STATE_REG_44,FROM_STATE_REG_45,FROM_STATE_REG_46,FROM_STATE_REG_47,FROM_STATE_REG_48,FROM_STATE_REG_49,FROM_STATE_REG_50,FROM_STATE_REG_51,FROM_STATE_REG_52,FROM_STATE_REG_53,FROM_STATE_REG_54,FROM_STATE_REG_55,FROM_STATE_REG_56,FROM_STATE_REG_57,FROM_STATE_REG_58,FROM_STATE_REG_59,FROM_STATE_REG_60,FROM_STATE_REG_61,FROM_STATE_REG_62,FROM_STATE_REG_63,FROM_STATE_REG_64,FROM_STATE_REG_65,FROM_STATE_REG_66,FROM_STATE_REG_67,FROM_STATE_REG_68,FROM_STATE_REG_69,FROM_STATE_REG_70,FROM_STATE_REG_71,FROM_STATE_REG_72,FROM_STATE_REG_73,FROM_STATE_REG_74,FROM_STATE_REG_75,FROM_STATE_REG_76,FROM_STATE_REG_77,FROM_STATE_REG_78,FROM_STATE_REG_79,FROM_STATE_REG_80,FROM_STATE_REG_81,FROM_STATE_REG_82,FROM_STATE_REG_83,FROM_STATE_REG_84,FROM_STATE_REG_85,FROM_STATE_REG_86,FROM_STATE_REG_87,FROM_STATE_REG_88,FROM_STATE_REG_89,FROM_STATE_REG_90,FROM_STATE_REG_91,FROM_STATE_REG_92,FROM_STATE_REG_93,FROM_STATE_REG_94,FROM_STATE_REG_95,FROM_STATE_REG_96,FROM_STATE_REG_97,FROM_STATE_REG_98,FROM_STATE_REG_99,FROM_STATE_REG_100,FROM_STATE_REG_101,FROM_STATE_REG_102,FROM_STATE_REG_103,FROM_STATE_REG_104,FROM_STATE_REG_105,FROM_STATE_REG_106,FROM_STATE_REG_107,FROM_STATE_REG_108,FROM_STATE_REG_109,FROM_STATE_REG_110,FROM_STATE_REG_111,FROM_STATE_REG_112,FROM_STATE_REG_113,FROM_STATE_REG_114,FROM_STATE_REG_115,FROM_STATE_REG_116,FROM_STATE_REG_117,FROM_STATE_REG_118,FROM_STATE_REG_119,FROM_STATE_REG_120,FROM_STATE_REG_121,FROM_STATE_REG_122,FROM_STATE_REG_123,FROM_STATE_REG_124,FROM_STATE_REG_125,FROM_STATE_REG_126,FROM_STATE_REG_127: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_SELECTION_UNIT_0,FROM_SELECTION_UNIT_1,FROM_SELECTION_UNIT_2,FROM_SELECTION_UNIT_3,FROM_SELECTION_UNIT_4,FROM_SELECTION_UNIT_5,FROM_SELECTION_UNIT_6,FROM_SELECTION_UNIT_7,FROM_SELECTION_UNIT_8,FROM_SELECTION_UNIT_9,FROM_SELECTION_UNIT_10,FROM_SELECTION_UNIT_11,FROM_SELECTION_UNIT_12,FROM_SELECTION_UNIT_13,FROM_SELECTION_UNIT_14,FROM_SELECTION_UNIT_15,FROM_SELECTION_UNIT_16,FROM_SELECTION_UNIT_17,FROM_SELECTION_UNIT_18,FROM_SELECTION_UNIT_19,FROM_SELECTION_UNIT_20,FROM_SELECTION_UNIT_21,FROM_SELECTION_UNIT_22,FROM_SELECTION_UNIT_23,FROM_SELECTION_UNIT_24,FROM_SELECTION_UNIT_25,FROM_SELECTION_UNIT_26,FROM_SELECTION_UNIT_27,FROM_SELECTION_UNIT_28,FROM_SELECTION_UNIT_29,FROM_SELECTION_UNIT_30,FROM_SELECTION_UNIT_31,FROM_SELECTION_UNIT_32,FROM_SELECTION_UNIT_33,FROM_SELECTION_UNIT_34,FROM_SELECTION_UNIT_35,FROM_SELECTION_UNIT_36,FROM_SELECTION_UNIT_37,FROM_SELECTION_UNIT_38,FROM_SELECTION_UNIT_39,FROM_SELECTION_UNIT_40,FROM_SELECTION_UNIT_41,FROM_SELECTION_UNIT_42,FROM_SELECTION_UNIT_43,FROM_SELECTION_UNIT_44,FROM_SELECTION_UNIT_45,FROM_SELECTION_UNIT_46,FROM_SELECTION_UNIT_47,FROM_SELECTION_UNIT_48,FROM_SELECTION_UNIT_49,FROM_SELECTION_UNIT_50,FROM_SELECTION_UNIT_51,FROM_SELECTION_UNIT_52,FROM_SELECTION_UNIT_53,FROM_SELECTION_UNIT_54,FROM_SELECTION_UNIT_55,FROM_SELECTION_UNIT_56,FROM_SELECTION_UNIT_57,FROM_SELECTION_UNIT_58,FROM_SELECTION_UNIT_59,FROM_SELECTION_UNIT_60,FROM_SELECTION_UNIT_61,FROM_SELECTION_UNIT_62,FROM_SELECTION_UNIT_63,FROM_SELECTION_UNIT_64,FROM_SELECTION_UNIT_65,FROM_SELECTION_UNIT_66,FROM_SELECTION_UNIT_67,FROM_SELECTION_UNIT_68,FROM_SELECTION_UNIT_69,FROM_SELECTION_UNIT_70,FROM_SELECTION_UNIT_71,FROM_SELECTION_UNIT_72,FROM_SELECTION_UNIT_73,FROM_SELECTION_UNIT_74,FROM_SELECTION_UNIT_75,FROM_SELECTION_UNIT_76,FROM_SELECTION_UNIT_77,FROM_SELECTION_UNIT_78,FROM_SELECTION_UNIT_79,FROM_SELECTION_UNIT_80,FROM_SELECTION_UNIT_81,FROM_SELECTION_UNIT_82,FROM_SELECTION_UNIT_83,FROM_SELECTION_UNIT_84,FROM_SELECTION_UNIT_85,FROM_SELECTION_UNIT_86,FROM_SELECTION_UNIT_87,FROM_SELECTION_UNIT_88,FROM_SELECTION_UNIT_89,FROM_SELECTION_UNIT_90,FROM_SELECTION_UNIT_91,FROM_SELECTION_UNIT_92,FROM_SELECTION_UNIT_93,FROM_SELECTION_UNIT_94,FROM_SELECTION_UNIT_95,FROM_SELECTION_UNIT_96,FROM_SELECTION_UNIT_97,FROM_SELECTION_UNIT_98,FROM_SELECTION_UNIT_99,FROM_SELECTION_UNIT_100,FROM_SELECTION_UNIT_101,FROM_SELECTION_UNIT_102,FROM_SELECTION_UNIT_103,FROM_SELECTION_UNIT_104,FROM_SELECTION_UNIT_105,FROM_SELECTION_UNIT_106,FROM_SELECTION_UNIT_107,FROM_SELECTION_UNIT_108,FROM_SELECTION_UNIT_109,FROM_SELECTION_UNIT_110,FROM_SELECTION_UNIT_111,FROM_SELECTION_UNIT_112,FROM_SELECTION_UNIT_113,FROM_SELECTION_UNIT_114,FROM_SELECTION_UNIT_115,FROM_SELECTION_UNIT_116,FROM_SELECTION_UNIT_117,FROM_SELECTION_UNIT_118,FROM_SELECTION_UNIT_119,FROM_SELECTION_UNIT_120,FROM_SELECTION_UNIT_121,FROM_SELECTION_UNIT_122,FROM_SELECTION_UNIT_123,FROM_SELECTION_UNIT_124,FROM_SELECTION_UNIT_125,FROM_SELECTION_UNIT_126,FROM_SELECTION_UNIT_127: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_0,FROM_WINDOW_1,FROM_WINDOW_2,FROM_WINDOW_3: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL MASKED_INPUT_0,MASKED_INPUT_2: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_DATAPATHS_0,FROM_DATAPATHS_1,FROM_DATAPATHS_2,FROM_DATAPATHS_3: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_CONTROL_UNITS_0,FROM_CONTROL_UNITS_1,FROM_CONTROL_UNITS_2,FROM_CONTROL_UNITS_3: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL UNWINDOWED_0,UNWINDOWED_1,UNWINDOWED_2,UNWINDOWED_3,UNWINDOWED_4,UNWINDOWED_5,UNWINDOWED_6,UNWINDOWED_7,UNWINDOWED_8,UNWINDOWED_9,UNWINDOWED_10,UNWINDOWED_11,UNWINDOWED_12,UNWINDOWED_13,UNWINDOWED_14,UNWINDOWED_15,UNWINDOWED_16,UNWINDOWED_17,UNWINDOWED_18,UNWINDOWED_19,UNWINDOWED_20,UNWINDOWED_21,UNWINDOWED_22,UNWINDOWED_23,UNWINDOWED_24,UNWINDOWED_25,UNWINDOWED_26,UNWINDOWED_27,UNWINDOWED_28,UNWINDOWED_29,UNWINDOWED_30,UNWINDOWED_31,UNWINDOWED_32,UNWINDOWED_33,UNWINDOWED_34,UNWINDOWED_35,UNWINDOWED_36,UNWINDOWED_37,UNWINDOWED_38,UNWINDOWED_39,UNWINDOWED_40,UNWINDOWED_41,UNWINDOWED_42,UNWINDOWED_43,UNWINDOWED_44,UNWINDOWED_45,UNWINDOWED_46,UNWINDOWED_47,UNWINDOWED_48,UNWINDOWED_49,UNWINDOWED_50,UNWINDOWED_51,UNWINDOWED_52,UNWINDOWED_53,UNWINDOWED_54,UNWINDOWED_55,UNWINDOWED_56,UNWINDOWED_57,UNWINDOWED_58,UNWINDOWED_59,UNWINDOWED_60,UNWINDOWED_61,UNWINDOWED_62,UNWINDOWED_63,UNWINDOWED_64,UNWINDOWED_65,UNWINDOWED_66,UNWINDOWED_67,UNWINDOWED_68,UNWINDOWED_69,UNWINDOWED_70,UNWINDOWED_71,UNWINDOWED_72,UNWINDOWED_73,UNWINDOWED_74,UNWINDOWED_75,UNWINDOWED_76,UNWINDOWED_77,UNWINDOWED_78,UNWINDOWED_79,UNWINDOWED_80,UNWINDOWED_81,UNWINDOWED_82,UNWINDOWED_83,UNWINDOWED_84,UNWINDOWED_85,UNWINDOWED_86,UNWINDOWED_87,UNWINDOWED_88,UNWINDOWED_89,UNWINDOWED_90,UNWINDOWED_91,UNWINDOWED_92,UNWINDOWED_93,UNWINDOWED_94,UNWINDOWED_95,UNWINDOWED_96,UNWINDOWED_97,UNWINDOWED_98,UNWINDOWED_99,UNWINDOWED_100,UNWINDOWED_101,UNWINDOWED_102,UNWINDOWED_103,UNWINDOWED_104,UNWINDOWED_105,UNWINDOWED_106,UNWINDOWED_107,UNWINDOWED_108,UNWINDOWED_109,UNWINDOWED_110,UNWINDOWED_111,UNWINDOWED_112,UNWINDOWED_113,UNWINDOWED_114,UNWINDOWED_115,UNWINDOWED_116,UNWINDOWED_117,UNWINDOWED_118,UNWINDOWED_119,UNWINDOWED_120,UNWINDOWED_121,UNWINDOWED_122,UNWINDOWED_123,UNWINDOWED_124,UNWINDOWED_125,UNWINDOWED_126,UNWINDOWED_127: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_DEC_MASK : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL UNWINDOWED_MASK, REORDERED_MASK, STATE_UPDATE_MASK : STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL SELECTED_OUTPUT: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_FIRST_CU_DONE : STD_LOGIC;

BEGIN

STATE_REG_0 : n_bit_register_clear_1
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_0 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(0) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_0);
STATE_REG_1 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1);
STATE_REG_2 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_2 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(2) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_2);
STATE_REG_3 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_3 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(3) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_3);
STATE_REG_4 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_4 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(4) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_4);
STATE_REG_5 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_5 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(5) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_5);
STATE_REG_6 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_6 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(6) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_6);
STATE_REG_7 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_7 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(7) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_7);
STATE_REG_8 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_8 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(8) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_8);
STATE_REG_9 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_9 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(9) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_9);
STATE_REG_10 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_10 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(10) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_10);
STATE_REG_11 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_11 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(11) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_11);
STATE_REG_12 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_12 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(12) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_12);
STATE_REG_13 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_13 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(13) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_13);
STATE_REG_14 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_14 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(14) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_14);
STATE_REG_15 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_15 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(15) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_15);
STATE_REG_16 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_16 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(16) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_16);
STATE_REG_17 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_17 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(17) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_17);
STATE_REG_18 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_18 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(18) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_18);
STATE_REG_19 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_19 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(19) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_19);
STATE_REG_20 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_20 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(20) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_20);
STATE_REG_21 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_21 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(21) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_21);
STATE_REG_22 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_22 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(22) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_22);
STATE_REG_23 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_23 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(23) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_23);
STATE_REG_24 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_24 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(24) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_24);
STATE_REG_25 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_25 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(25) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_25);
STATE_REG_26 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_26 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(26) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_26);
STATE_REG_27 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_27 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(27) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_27);
STATE_REG_28 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_28 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(28) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_28);
STATE_REG_29 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_29 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(29) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_29);
STATE_REG_30 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_30 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(30) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_30);
STATE_REG_31 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_31 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(31) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_31);
STATE_REG_32 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_32 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(32) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_32);
STATE_REG_33 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_33 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(33) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_33);
STATE_REG_34 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_34 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(34) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_34);
STATE_REG_35 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_35 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(35) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_35);
STATE_REG_36 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_36 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(36) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_36);
STATE_REG_37 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_37 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(37) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_37);
STATE_REG_38 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_38 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(38) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_38);
STATE_REG_39 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_39 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(39) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_39);
STATE_REG_40 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_40 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(40) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_40);
STATE_REG_41 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_41 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(41) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_41);
STATE_REG_42 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_42 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(42) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_42);
STATE_REG_43 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_43 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(43) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_43);
STATE_REG_44 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_44 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(44) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_44);
STATE_REG_45 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_45 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(45) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_45);
STATE_REG_46 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_46 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(46) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_46);
STATE_REG_47 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_47 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(47) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_47);
STATE_REG_48 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_48 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(48) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_48);
STATE_REG_49 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_49 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(49) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_49);
STATE_REG_50 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_50 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(50) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_50);
STATE_REG_51 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_51 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(51) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_51);
STATE_REG_52 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_52 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(52) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_52);
STATE_REG_53 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_53 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(53) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_53);
STATE_REG_54 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_54 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(54) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_54);
STATE_REG_55 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_55 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(55) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_55);
STATE_REG_56 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_56 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(56) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_56);
STATE_REG_57 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_57 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(57) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_57);
STATE_REG_58 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_58 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(58) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_58);
STATE_REG_59 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_59 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(59) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_59);
STATE_REG_60 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_60 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(60) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_60);
STATE_REG_61 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_61 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(61) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_61);
STATE_REG_62 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_62 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(62) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_62);
STATE_REG_63 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_63 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(63) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_63);
STATE_REG_64 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_64 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(64) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_64);
STATE_REG_65 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_65 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(65) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_65);
STATE_REG_66 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_66 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(66) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_66);
STATE_REG_67 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_67 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(67) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_67);
STATE_REG_68 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_68 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(68) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_68);
STATE_REG_69 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_69 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(69) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_69);
STATE_REG_70 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_70 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(70) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_70);
STATE_REG_71 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_71 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(71) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_71);
STATE_REG_72 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_72 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(72) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_72);
STATE_REG_73 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_73 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(73) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_73);
STATE_REG_74 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_74 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(74) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_74);
STATE_REG_75 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_75 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(75) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_75);
STATE_REG_76 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_76 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(76) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_76);
STATE_REG_77 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_77 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(77) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_77);
STATE_REG_78 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_78 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(78) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_78);
STATE_REG_79 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_79 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(79) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_79);
STATE_REG_80 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_80 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(80) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_80);
STATE_REG_81 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_81 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(81) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_81);
STATE_REG_82 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_82 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(82) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_82);
STATE_REG_83 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_83 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(83) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_83);
STATE_REG_84 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_84 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(84) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_84);
STATE_REG_85 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_85 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(85) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_85);
STATE_REG_86 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_86 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(86) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_86);
STATE_REG_87 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_87 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(87) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_87);
STATE_REG_88 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_88 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(88) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_88);
STATE_REG_89 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_89 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(89) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_89);
STATE_REG_90 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_90 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(90) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_90);
STATE_REG_91 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_91 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(91) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_91);
STATE_REG_92 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_92 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(92) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_92);
STATE_REG_93 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_93 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(93) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_93);
STATE_REG_94 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_94 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(94) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_94);
STATE_REG_95 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_95 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(95) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_95);
STATE_REG_96 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_96 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(96) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_96);
STATE_REG_97 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_97 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(97) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_97);
STATE_REG_98 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_98 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(98) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_98);
STATE_REG_99 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_99 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(99) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_99);
STATE_REG_100 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_100 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(100) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_100);
STATE_REG_101 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_101 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(101) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_101);
STATE_REG_102 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_102 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(102) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_102);
STATE_REG_103 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_103 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(103) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_103);
STATE_REG_104 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_104 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(104) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_104);
STATE_REG_105 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_105 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(105) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_105);
STATE_REG_106 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_106 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(106) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_106);
STATE_REG_107 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_107 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(107) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_107);
STATE_REG_108 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_108 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(108) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_108);
STATE_REG_109 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_109 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(109) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_109);
STATE_REG_110 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_110 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(110) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_110);
STATE_REG_111 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_111 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(111) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_111);
STATE_REG_112 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_112 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(112) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_112);
STATE_REG_113 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_113 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(113) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_113);
STATE_REG_114 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_114 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(114) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_114);
STATE_REG_115 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_115 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(115) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_115);
STATE_REG_116 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_116 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(116) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_116);
STATE_REG_117 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_117 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(117) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_117);
STATE_REG_118 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_118 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(118) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_118);
STATE_REG_119 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_119 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(119) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_119);
STATE_REG_120 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_120 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(120) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_120);
STATE_REG_121 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_121 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(121) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_121);
STATE_REG_122 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_122 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(122) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_122);
STATE_REG_123 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_123 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(123) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_123);
STATE_REG_124 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_124 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(124) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_124);
STATE_REG_125 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_125 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(125) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_125);
STATE_REG_126 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_126 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(126) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_126);
STATE_REG_127 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_127 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(127) ,
												REG_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_127);


MUX_SEL_UNIT_0 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_0 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_0 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_0 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_0 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_0 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_0 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_0
									);
MUX_SEL_UNIT_1 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_1 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_2 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_4 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_8 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_16 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_32 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_64 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_1
									);
MUX_SEL_UNIT_2 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_2 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_1 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_1 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_1 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_1 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_1 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_2
									);
MUX_SEL_UNIT_3 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_3 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_3 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_5 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_9 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_17 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_33 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_65 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_3
									);
MUX_SEL_UNIT_4 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_4 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_4 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_2 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_2 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_2 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_2 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_4
									);
MUX_SEL_UNIT_5 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_5 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_6 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_6 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_10 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_18 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_34 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_66 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_5
									);
MUX_SEL_UNIT_6 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_6 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_5 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_3 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_3 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_3 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_3 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_6
									);
MUX_SEL_UNIT_7 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_7 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_7 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_7 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_11 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_19 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_35 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_67 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_7
									);
MUX_SEL_UNIT_8 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_8 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_8 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_8 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_4 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_4 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_4 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_8
									);
MUX_SEL_UNIT_9 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_9 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_10 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_12 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_12 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_20 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_36 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_68 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_9
									);
MUX_SEL_UNIT_10 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_10 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_9 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_9 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_5 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_5 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_5 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_5 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_10
									);
MUX_SEL_UNIT_11 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_11 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_11 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_13 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_13 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_21 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_37 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_69 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_11
									);
MUX_SEL_UNIT_12 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_12 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_12 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_10 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_6 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_6 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_6 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_6 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_12
									);
MUX_SEL_UNIT_13 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_13 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_14 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_14 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_14 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_22 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_38 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_70 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_13
									);
MUX_SEL_UNIT_14 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_14 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_13 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_11 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_7 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_7 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_7 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_7 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_14
									);
MUX_SEL_UNIT_15 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_15 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_15 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_15 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_15 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_23 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_39 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_71 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_15
									);
MUX_SEL_UNIT_16 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_16 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_16 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_16 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_16 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_8 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_8 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_8 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_16
									);
MUX_SEL_UNIT_17 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_17 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_18 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_20 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_24 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_24 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_40 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_72 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_17
									);
MUX_SEL_UNIT_18 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_18 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_17 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_17 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_17 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_9 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_9 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_9 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_18
									);
MUX_SEL_UNIT_19 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_19 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_19 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_21 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_25 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_25 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_41 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_73 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_19
									);
MUX_SEL_UNIT_20 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_20 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_20 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_18 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_18 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_10 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_10 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_10 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_20
									);
MUX_SEL_UNIT_21 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_21 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_22 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_22 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_26 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_26 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_42 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_74 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_21
									);
MUX_SEL_UNIT_22 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_22 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_21 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_19 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_19 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_11 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_11 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_11 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_22
									);
MUX_SEL_UNIT_23 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_23 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_23 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_23 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_27 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_27 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_43 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_75 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_23
									);
MUX_SEL_UNIT_24 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_24 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_24 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_24 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_20 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_12 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_12 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_12 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_24
									);
MUX_SEL_UNIT_25 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_25 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_26 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_28 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_28 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_28 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_44 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_76 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_25
									);
MUX_SEL_UNIT_26 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_26 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_25 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_25 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_21 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_13 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_13 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_13 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_26
									);
MUX_SEL_UNIT_27 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_27 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_27 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_29 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_29 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_29 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_45 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_77 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_27
									);
MUX_SEL_UNIT_28 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_28 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_28 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_26 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_22 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_14 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_14 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_14 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_28
									);
MUX_SEL_UNIT_29 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_29 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_30 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_30 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_30 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_30 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_46 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_78 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_29
									);
MUX_SEL_UNIT_30 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_30 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_29 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_27 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_23 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_15 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_15 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_15 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_30
									);
MUX_SEL_UNIT_31 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_31 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_31 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_31 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_31 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_31 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_47 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_79 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_31
									);
MUX_SEL_UNIT_32 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_32 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_32 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_32 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_32 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_32 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_16 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_16 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_32
									);
MUX_SEL_UNIT_33 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_33 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_34 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_36 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_40 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_48 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_48 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_80 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_33
									);
MUX_SEL_UNIT_34 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_34 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_33 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_33 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_33 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_33 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_17 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_17 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_34
									);
MUX_SEL_UNIT_35 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_35 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_35 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_37 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_41 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_49 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_49 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_81 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_35
									);
MUX_SEL_UNIT_36 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_36 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_36 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_34 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_34 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_34 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_18 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_18 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_36
									);
MUX_SEL_UNIT_37 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_37 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_38 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_38 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_42 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_50 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_50 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_82 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_37
									);
MUX_SEL_UNIT_38 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_38 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_37 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_35 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_35 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_35 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_19 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_19 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_38
									);
MUX_SEL_UNIT_39 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_39 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_39 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_39 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_43 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_51 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_51 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_83 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_39
									);
MUX_SEL_UNIT_40 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_40 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_40 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_40 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_36 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_36 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_20 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_20 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_40
									);
MUX_SEL_UNIT_41 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_41 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_42 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_44 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_44 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_52 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_52 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_84 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_41
									);
MUX_SEL_UNIT_42 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_42 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_41 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_41 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_37 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_37 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_21 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_21 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_42
									);
MUX_SEL_UNIT_43 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_43 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_43 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_45 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_45 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_53 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_53 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_85 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_43
									);
MUX_SEL_UNIT_44 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_44 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_44 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_42 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_38 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_38 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_22 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_22 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_44
									);
MUX_SEL_UNIT_45 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_45 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_46 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_46 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_46 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_54 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_54 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_86 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_45
									);
MUX_SEL_UNIT_46 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_46 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_45 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_43 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_39 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_39 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_23 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_23 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_46
									);
MUX_SEL_UNIT_47 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_47 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_47 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_47 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_47 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_55 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_55 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_87 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_47
									);
MUX_SEL_UNIT_48 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_48 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_48 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_48 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_48 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_40 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_24 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_24 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_48
									);
MUX_SEL_UNIT_49 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_49 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_50 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_52 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_56 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_56 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_56 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_88 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_49
									);
MUX_SEL_UNIT_50 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_50 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_49 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_49 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_49 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_41 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_25 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_25 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_50
									);
MUX_SEL_UNIT_51 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_51 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_51 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_53 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_57 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_57 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_57 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_89 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_51
									);
MUX_SEL_UNIT_52 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_52 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_52 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_50 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_50 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_42 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_26 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_26 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_52
									);
MUX_SEL_UNIT_53 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_53 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_54 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_54 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_58 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_58 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_58 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_90 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_53
									);
MUX_SEL_UNIT_54 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_54 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_53 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_51 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_51 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_43 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_27 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_27 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_54
									);
MUX_SEL_UNIT_55 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_55 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_55 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_55 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_59 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_59 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_59 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_91 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_55
									);
MUX_SEL_UNIT_56 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_56 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_56 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_56 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_52 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_44 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_28 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_28 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_56
									);
MUX_SEL_UNIT_57 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_57 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_58 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_60 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_60 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_60 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_60 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_92 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_57
									);
MUX_SEL_UNIT_58 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_58 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_57 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_57 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_53 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_45 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_29 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_29 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_58
									);
MUX_SEL_UNIT_59 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_59 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_59 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_61 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_61 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_61 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_61 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_93 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_59
									);
MUX_SEL_UNIT_60 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_60 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_60 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_58 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_54 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_46 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_30 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_30 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_60
									);
MUX_SEL_UNIT_61 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_61 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_62 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_62 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_62 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_62 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_62 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_94 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_61
									);
MUX_SEL_UNIT_62 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_62 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_61 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_59 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_55 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_47 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_31 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_31 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_62
									);
MUX_SEL_UNIT_63 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_63 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_63 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_63 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_63 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_63 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_63 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_95 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_63
									);
MUX_SEL_UNIT_64 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_64 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_64 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_64 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_64 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_64 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_64 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_32 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_64
									);
MUX_SEL_UNIT_65 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_65 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_66 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_68 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_72 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_80 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_96 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_96 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_65
									);
MUX_SEL_UNIT_66 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_66 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_65 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_65 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_65 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_65 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_65 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_33 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_66
									);
MUX_SEL_UNIT_67 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_67 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_67 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_69 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_73 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_81 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_97 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_97 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_67
									);
MUX_SEL_UNIT_68 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_68 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_68 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_66 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_66 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_66 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_66 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_34 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_68
									);
MUX_SEL_UNIT_69 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_69 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_70 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_70 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_74 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_82 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_98 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_98 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_69
									);
MUX_SEL_UNIT_70 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_70 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_69 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_67 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_67 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_67 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_67 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_35 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_70
									);
MUX_SEL_UNIT_71 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_71 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_71 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_71 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_75 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_83 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_99 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_99 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_71
									);
MUX_SEL_UNIT_72 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_72 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_72 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_72 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_68 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_68 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_68 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_36 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_72
									);
MUX_SEL_UNIT_73 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_73 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_74 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_76 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_76 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_84 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_100 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_100 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_73
									);
MUX_SEL_UNIT_74 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_74 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_73 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_73 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_69 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_69 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_69 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_37 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_74
									);
MUX_SEL_UNIT_75 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_75 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_75 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_77 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_77 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_85 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_101 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_101 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_75
									);
MUX_SEL_UNIT_76 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_76 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_76 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_74 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_70 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_70 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_70 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_38 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_76
									);
MUX_SEL_UNIT_77 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_77 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_78 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_78 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_78 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_86 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_102 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_102 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_77
									);
MUX_SEL_UNIT_78 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_78 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_77 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_75 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_71 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_71 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_71 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_39 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_78
									);
MUX_SEL_UNIT_79 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_79 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_79 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_79 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_79 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_87 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_103 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_103 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_79
									);
MUX_SEL_UNIT_80 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_80 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_80 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_80 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_80 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_72 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_72 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_40 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_80
									);
MUX_SEL_UNIT_81 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_81 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_82 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_84 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_88 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_88 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_104 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_104 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_81
									);
MUX_SEL_UNIT_82 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_82 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_81 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_81 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_81 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_73 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_73 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_41 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_82
									);
MUX_SEL_UNIT_83 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_83 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_83 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_85 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_89 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_89 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_105 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_105 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_83
									);
MUX_SEL_UNIT_84 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_84 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_84 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_82 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_82 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_74 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_74 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_42 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_84
									);
MUX_SEL_UNIT_85 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_85 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_86 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_86 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_90 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_90 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_106 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_106 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_85
									);
MUX_SEL_UNIT_86 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_86 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_85 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_83 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_83 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_75 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_75 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_43 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_86
									);
MUX_SEL_UNIT_87 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_87 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_87 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_87 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_91 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_91 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_107 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_107 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_87
									);
MUX_SEL_UNIT_88 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_88 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_88 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_88 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_84 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_76 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_76 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_44 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_88
									);
MUX_SEL_UNIT_89 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_89 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_90 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_92 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_92 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_92 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_108 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_108 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_89
									);
MUX_SEL_UNIT_90 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_90 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_89 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_89 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_85 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_77 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_77 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_45 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_90
									);
MUX_SEL_UNIT_91 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_91 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_91 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_93 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_93 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_93 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_109 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_109 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_91
									);
MUX_SEL_UNIT_92 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_92 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_92 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_90 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_86 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_78 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_78 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_46 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_92
									);
MUX_SEL_UNIT_93 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_93 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_94 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_94 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_94 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_94 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_110 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_110 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_93
									);
MUX_SEL_UNIT_94 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_94 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_93 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_91 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_87 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_79 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_79 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_47 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_94
									);
MUX_SEL_UNIT_95 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_95 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_95 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_95 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_95 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_95 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_111 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_111 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_95
									);
MUX_SEL_UNIT_96 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_96 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_96 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_96 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_96 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_96 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_80 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_48 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_96
									);
MUX_SEL_UNIT_97 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_97 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_98 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_100 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_104 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_112 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_112 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_112 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_97
									);
MUX_SEL_UNIT_98 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_98 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_97 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_97 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_97 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_97 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_81 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_49 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_98
									);
MUX_SEL_UNIT_99 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_99 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_99 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_101 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_105 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_113 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_113 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_113 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_99
									);
MUX_SEL_UNIT_100 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_100 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_100 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_98 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_98 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_98 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_82 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_50 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_100
									);
MUX_SEL_UNIT_101 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_101 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_102 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_102 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_106 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_114 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_114 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_114 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_101
									);
MUX_SEL_UNIT_102 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_102 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_101 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_99 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_99 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_99 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_83 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_51 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_102
									);
MUX_SEL_UNIT_103 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_103 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_103 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_103 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_107 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_115 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_115 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_115 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_103
									);
MUX_SEL_UNIT_104 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_104 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_104 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_104 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_100 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_100 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_84 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_52 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_104
									);
MUX_SEL_UNIT_105 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_105 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_106 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_108 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_108 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_116 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_116 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_116 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_105
									);
MUX_SEL_UNIT_106 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_106 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_105 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_105 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_101 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_101 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_85 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_53 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_106
									);
MUX_SEL_UNIT_107 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_107 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_107 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_109 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_109 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_117 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_117 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_117 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_107
									);
MUX_SEL_UNIT_108 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_108 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_108 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_106 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_102 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_102 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_86 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_54 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_108
									);
MUX_SEL_UNIT_109 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_109 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_110 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_110 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_110 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_118 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_118 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_118 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_109
									);
MUX_SEL_UNIT_110 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_110 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_109 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_107 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_103 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_103 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_87 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_55 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_110
									);
MUX_SEL_UNIT_111 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_111 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_111 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_111 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_111 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_119 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_119 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_119 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_111
									);
MUX_SEL_UNIT_112 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_112 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_112 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_112 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_112 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_104 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_88 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_56 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_112
									);
MUX_SEL_UNIT_113 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_113 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_114 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_116 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_120 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_120 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_120 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_120 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_113
									);
MUX_SEL_UNIT_114 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_114 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_113 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_113 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_113 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_105 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_89 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_57 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_114
									);
MUX_SEL_UNIT_115 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_115 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_115 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_117 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_121 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_121 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_121 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_121 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_115
									);
MUX_SEL_UNIT_116 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_116 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_116 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_114 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_114 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_106 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_90 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_58 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_116
									);
MUX_SEL_UNIT_117 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_117 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_118 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_118 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_122 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_122 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_122 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_122 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_117
									);
MUX_SEL_UNIT_118 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_118 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_117 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_115 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_115 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_107 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_91 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_59 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_118
									);
MUX_SEL_UNIT_119 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_119 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_119 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_119 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_123 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_123 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_123 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_123 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_119
									);
MUX_SEL_UNIT_120 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_120 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_120 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_120 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_116 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_108 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_92 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_60 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_120
									);
MUX_SEL_UNIT_121 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_121 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_122 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_124 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_124 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_124 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_124 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_124 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_121
									);
MUX_SEL_UNIT_122 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_122 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_121 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_121 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_117 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_109 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_93 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_61 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_122
									);
MUX_SEL_UNIT_123 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_123 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_123 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_125 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_125 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_125 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_125 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_125 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_123
									);
MUX_SEL_UNIT_124 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_124 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_124 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_122 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_118 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_110 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_94 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_62 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_124
									);
MUX_SEL_UNIT_125 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_125 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_126 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_126 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_126 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_126 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_126 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_126 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_125
									);
MUX_SEL_UNIT_126 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_126 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_125 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_123 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_119 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_111 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_95 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_63 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_126
									);
MUX_SEL_UNIT_127 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => FROM_STATE_REG_127 ,
										MUX_7_1_IN_1 => FROM_STATE_REG_127 ,
										MUX_7_1_IN_2 => FROM_STATE_REG_127 ,
										MUX_7_1_IN_3 => FROM_STATE_REG_127 ,
										MUX_7_1_IN_4 => FROM_STATE_REG_127 ,
										MUX_7_1_IN_5 => FROM_STATE_REG_127 ,
										MUX_7_1_IN_6 => FROM_STATE_REG_127 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => FROM_SELECTION_UNIT_127
									);

MUX_WINDOWING_UNIT_0 : multiplexer_32_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_32_1_IN_0 => FROM_SELECTION_UNIT_0 ,
										MUX_32_1_IN_1 => FROM_SELECTION_UNIT_4 ,
										MUX_32_1_IN_2 => FROM_SELECTION_UNIT_8 ,
										MUX_32_1_IN_3 => FROM_SELECTION_UNIT_12 ,
										MUX_32_1_IN_4 => FROM_SELECTION_UNIT_16 ,
										MUX_32_1_IN_5 => FROM_SELECTION_UNIT_20 ,
										MUX_32_1_IN_6 => FROM_SELECTION_UNIT_24 ,
										MUX_32_1_IN_7 => FROM_SELECTION_UNIT_28 ,
										MUX_32_1_IN_8 => FROM_SELECTION_UNIT_32 ,
										MUX_32_1_IN_9 => FROM_SELECTION_UNIT_36 ,
										MUX_32_1_IN_10 => FROM_SELECTION_UNIT_40 ,
										MUX_32_1_IN_11 => FROM_SELECTION_UNIT_44 ,
										MUX_32_1_IN_12 => FROM_SELECTION_UNIT_48 ,
										MUX_32_1_IN_13 => FROM_SELECTION_UNIT_52 ,
										MUX_32_1_IN_14 => FROM_SELECTION_UNIT_56 ,
										MUX_32_1_IN_15 => FROM_SELECTION_UNIT_60 ,
										MUX_32_1_IN_16 => FROM_SELECTION_UNIT_64 ,
										MUX_32_1_IN_17 => FROM_SELECTION_UNIT_68 ,
										MUX_32_1_IN_18 => FROM_SELECTION_UNIT_72 ,
										MUX_32_1_IN_19 => FROM_SELECTION_UNIT_76 ,
										MUX_32_1_IN_20 => FROM_SELECTION_UNIT_80 ,
										MUX_32_1_IN_21 => FROM_SELECTION_UNIT_84 ,
										MUX_32_1_IN_22 => FROM_SELECTION_UNIT_88 ,
										MUX_32_1_IN_23 => FROM_SELECTION_UNIT_92 ,
										MUX_32_1_IN_24 => FROM_SELECTION_UNIT_96 ,
										MUX_32_1_IN_25 => FROM_SELECTION_UNIT_100 ,
										MUX_32_1_IN_26 => FROM_SELECTION_UNIT_104 ,
										MUX_32_1_IN_27 => FROM_SELECTION_UNIT_108 ,
										MUX_32_1_IN_28 => FROM_SELECTION_UNIT_112 ,
										MUX_32_1_IN_29 => FROM_SELECTION_UNIT_116 ,
										MUX_32_1_IN_30 => FROM_SELECTION_UNIT_120 ,
										MUX_32_1_IN_31 => FROM_SELECTION_UNIT_124 ,
				                    			MUX_32_1_IN_SEL => QEP_N_7_W_5_S_0_IN_WIN_SEL ,
										MUX_32_1_OUT_RES => FROM_WINDOW_0
									);
MUX_WINDOWING_UNIT_1 : multiplexer_32_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_32_1_IN_0 => FROM_SELECTION_UNIT_1 ,
										MUX_32_1_IN_1 => FROM_SELECTION_UNIT_5 ,
										MUX_32_1_IN_2 => FROM_SELECTION_UNIT_9 ,
										MUX_32_1_IN_3 => FROM_SELECTION_UNIT_13 ,
										MUX_32_1_IN_4 => FROM_SELECTION_UNIT_17 ,
										MUX_32_1_IN_5 => FROM_SELECTION_UNIT_21 ,
										MUX_32_1_IN_6 => FROM_SELECTION_UNIT_25 ,
										MUX_32_1_IN_7 => FROM_SELECTION_UNIT_29 ,
										MUX_32_1_IN_8 => FROM_SELECTION_UNIT_33 ,
										MUX_32_1_IN_9 => FROM_SELECTION_UNIT_37 ,
										MUX_32_1_IN_10 => FROM_SELECTION_UNIT_41 ,
										MUX_32_1_IN_11 => FROM_SELECTION_UNIT_45 ,
										MUX_32_1_IN_12 => FROM_SELECTION_UNIT_49 ,
										MUX_32_1_IN_13 => FROM_SELECTION_UNIT_53 ,
										MUX_32_1_IN_14 => FROM_SELECTION_UNIT_57 ,
										MUX_32_1_IN_15 => FROM_SELECTION_UNIT_61 ,
										MUX_32_1_IN_16 => FROM_SELECTION_UNIT_65 ,
										MUX_32_1_IN_17 => FROM_SELECTION_UNIT_69 ,
										MUX_32_1_IN_18 => FROM_SELECTION_UNIT_73 ,
										MUX_32_1_IN_19 => FROM_SELECTION_UNIT_77 ,
										MUX_32_1_IN_20 => FROM_SELECTION_UNIT_81 ,
										MUX_32_1_IN_21 => FROM_SELECTION_UNIT_85 ,
										MUX_32_1_IN_22 => FROM_SELECTION_UNIT_89 ,
										MUX_32_1_IN_23 => FROM_SELECTION_UNIT_93 ,
										MUX_32_1_IN_24 => FROM_SELECTION_UNIT_97 ,
										MUX_32_1_IN_25 => FROM_SELECTION_UNIT_101 ,
										MUX_32_1_IN_26 => FROM_SELECTION_UNIT_105 ,
										MUX_32_1_IN_27 => FROM_SELECTION_UNIT_109 ,
										MUX_32_1_IN_28 => FROM_SELECTION_UNIT_113 ,
										MUX_32_1_IN_29 => FROM_SELECTION_UNIT_117 ,
										MUX_32_1_IN_30 => FROM_SELECTION_UNIT_121 ,
										MUX_32_1_IN_31 => FROM_SELECTION_UNIT_125 ,
				                    			MUX_32_1_IN_SEL => QEP_N_7_W_5_S_0_IN_WIN_SEL ,
										MUX_32_1_OUT_RES => FROM_WINDOW_1
									);
MUX_WINDOWING_UNIT_2 : multiplexer_32_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_32_1_IN_0 => FROM_SELECTION_UNIT_2 ,
										MUX_32_1_IN_1 => FROM_SELECTION_UNIT_6 ,
										MUX_32_1_IN_2 => FROM_SELECTION_UNIT_10 ,
										MUX_32_1_IN_3 => FROM_SELECTION_UNIT_14 ,
										MUX_32_1_IN_4 => FROM_SELECTION_UNIT_18 ,
										MUX_32_1_IN_5 => FROM_SELECTION_UNIT_22 ,
										MUX_32_1_IN_6 => FROM_SELECTION_UNIT_26 ,
										MUX_32_1_IN_7 => FROM_SELECTION_UNIT_30 ,
										MUX_32_1_IN_8 => FROM_SELECTION_UNIT_34 ,
										MUX_32_1_IN_9 => FROM_SELECTION_UNIT_38 ,
										MUX_32_1_IN_10 => FROM_SELECTION_UNIT_42 ,
										MUX_32_1_IN_11 => FROM_SELECTION_UNIT_46 ,
										MUX_32_1_IN_12 => FROM_SELECTION_UNIT_50 ,
										MUX_32_1_IN_13 => FROM_SELECTION_UNIT_54 ,
										MUX_32_1_IN_14 => FROM_SELECTION_UNIT_58 ,
										MUX_32_1_IN_15 => FROM_SELECTION_UNIT_62 ,
										MUX_32_1_IN_16 => FROM_SELECTION_UNIT_66 ,
										MUX_32_1_IN_17 => FROM_SELECTION_UNIT_70 ,
										MUX_32_1_IN_18 => FROM_SELECTION_UNIT_74 ,
										MUX_32_1_IN_19 => FROM_SELECTION_UNIT_78 ,
										MUX_32_1_IN_20 => FROM_SELECTION_UNIT_82 ,
										MUX_32_1_IN_21 => FROM_SELECTION_UNIT_86 ,
										MUX_32_1_IN_22 => FROM_SELECTION_UNIT_90 ,
										MUX_32_1_IN_23 => FROM_SELECTION_UNIT_94 ,
										MUX_32_1_IN_24 => FROM_SELECTION_UNIT_98 ,
										MUX_32_1_IN_25 => FROM_SELECTION_UNIT_102 ,
										MUX_32_1_IN_26 => FROM_SELECTION_UNIT_106 ,
										MUX_32_1_IN_27 => FROM_SELECTION_UNIT_110 ,
										MUX_32_1_IN_28 => FROM_SELECTION_UNIT_114 ,
										MUX_32_1_IN_29 => FROM_SELECTION_UNIT_118 ,
										MUX_32_1_IN_30 => FROM_SELECTION_UNIT_122 ,
										MUX_32_1_IN_31 => FROM_SELECTION_UNIT_126 ,
				                    			MUX_32_1_IN_SEL => QEP_N_7_W_5_S_0_IN_WIN_SEL ,
										MUX_32_1_OUT_RES => FROM_WINDOW_2
									);
MUX_WINDOWING_UNIT_3 : multiplexer_32_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_32_1_IN_0 => FROM_SELECTION_UNIT_3 ,
										MUX_32_1_IN_1 => FROM_SELECTION_UNIT_7 ,
										MUX_32_1_IN_2 => FROM_SELECTION_UNIT_11 ,
										MUX_32_1_IN_3 => FROM_SELECTION_UNIT_15 ,
										MUX_32_1_IN_4 => FROM_SELECTION_UNIT_19 ,
										MUX_32_1_IN_5 => FROM_SELECTION_UNIT_23 ,
										MUX_32_1_IN_6 => FROM_SELECTION_UNIT_27 ,
										MUX_32_1_IN_7 => FROM_SELECTION_UNIT_31 ,
										MUX_32_1_IN_8 => FROM_SELECTION_UNIT_35 ,
										MUX_32_1_IN_9 => FROM_SELECTION_UNIT_39 ,
										MUX_32_1_IN_10 => FROM_SELECTION_UNIT_43 ,
										MUX_32_1_IN_11 => FROM_SELECTION_UNIT_47 ,
										MUX_32_1_IN_12 => FROM_SELECTION_UNIT_51 ,
										MUX_32_1_IN_13 => FROM_SELECTION_UNIT_55 ,
										MUX_32_1_IN_14 => FROM_SELECTION_UNIT_59 ,
										MUX_32_1_IN_15 => FROM_SELECTION_UNIT_63 ,
										MUX_32_1_IN_16 => FROM_SELECTION_UNIT_67 ,
										MUX_32_1_IN_17 => FROM_SELECTION_UNIT_71 ,
										MUX_32_1_IN_18 => FROM_SELECTION_UNIT_75 ,
										MUX_32_1_IN_19 => FROM_SELECTION_UNIT_79 ,
										MUX_32_1_IN_20 => FROM_SELECTION_UNIT_83 ,
										MUX_32_1_IN_21 => FROM_SELECTION_UNIT_87 ,
										MUX_32_1_IN_22 => FROM_SELECTION_UNIT_91 ,
										MUX_32_1_IN_23 => FROM_SELECTION_UNIT_95 ,
										MUX_32_1_IN_24 => FROM_SELECTION_UNIT_99 ,
										MUX_32_1_IN_25 => FROM_SELECTION_UNIT_103 ,
										MUX_32_1_IN_26 => FROM_SELECTION_UNIT_107 ,
										MUX_32_1_IN_27 => FROM_SELECTION_UNIT_111 ,
										MUX_32_1_IN_28 => FROM_SELECTION_UNIT_115 ,
										MUX_32_1_IN_29 => FROM_SELECTION_UNIT_119 ,
										MUX_32_1_IN_30 => FROM_SELECTION_UNIT_123 ,
										MUX_32_1_IN_31 => FROM_SELECTION_UNIT_127 ,
				                    			MUX_32_1_IN_SEL => QEP_N_7_W_5_S_0_IN_WIN_SEL ,
										MUX_32_1_OUT_RES => FROM_WINDOW_3
									);
MASKED_INPUT_0 <= FROM_WINDOW_0 WHEN QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_2 <= FROM_WINDOW_2 WHEN QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');

FROM_WINDOW_DEC_MASK <= 
"00000000000000000000000000000001" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00000" ELSE
"00000000000000000000000000000010" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00001" ELSE
"00000000000000000000000000000100" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00010" ELSE
"00000000000000000000000000001000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00011" ELSE
"00000000000000000000000000010000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00100" ELSE
"00000000000000000000000000100000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00101" ELSE
"00000000000000000000000001000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00110" ELSE
"00000000000000000000000010000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "00111" ELSE
"00000000000000000000000100000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01000" ELSE
"00000000000000000000001000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01001" ELSE
"00000000000000000000010000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01010" ELSE
"00000000000000000000100000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01011" ELSE
"00000000000000000001000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01100" ELSE
"00000000000000000010000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01101" ELSE
"00000000000000000100000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01110" ELSE
"00000000000000001000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "01111" ELSE
"00000000000000010000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10000" ELSE
"00000000000000100000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10001" ELSE
"00000000000001000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10010" ELSE
"00000000000010000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10011" ELSE
"00000000000100000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10100" ELSE
"00000000001000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10101" ELSE
"00000000010000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10110" ELSE
"00000000100000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "10111" ELSE
"00000001000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11000" ELSE
"00000010000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11001" ELSE
"00000100000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11010" ELSE
"00001000000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11011" ELSE
"00010000000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11100" ELSE
"00100000000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11101" ELSE
"01000000000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11110" ELSE
"10000000000000000000000000000000" WHEN QEP_N_7_W_5_S_0_IN_WIN_SEL = "11111" ELSE
(OTHERS => '0');

UNWINDOWED_MASK(0) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(2) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(3) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(4) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(5) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(6) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(7) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(8) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(9) <= FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(10) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(11) <= FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(12) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(13) <= FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(14) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(15) <= FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(16) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(17) <= FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(18) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(19) <= FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(20) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(21) <= FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(22) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(23) <= FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(24) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(25) <= FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(26) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(27) <= FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(28) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(29) <= FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(30) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(31) <= FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(32) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(8);
UNWINDOWED_MASK(33) <= FROM_WINDOW_DEC_MASK(8);
UNWINDOWED_MASK(34) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(8);
UNWINDOWED_MASK(35) <= FROM_WINDOW_DEC_MASK(8);
UNWINDOWED_MASK(36) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(9);
UNWINDOWED_MASK(37) <= FROM_WINDOW_DEC_MASK(9);
UNWINDOWED_MASK(38) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(9);
UNWINDOWED_MASK(39) <= FROM_WINDOW_DEC_MASK(9);
UNWINDOWED_MASK(40) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(10);
UNWINDOWED_MASK(41) <= FROM_WINDOW_DEC_MASK(10);
UNWINDOWED_MASK(42) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(10);
UNWINDOWED_MASK(43) <= FROM_WINDOW_DEC_MASK(10);
UNWINDOWED_MASK(44) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(11);
UNWINDOWED_MASK(45) <= FROM_WINDOW_DEC_MASK(11);
UNWINDOWED_MASK(46) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(11);
UNWINDOWED_MASK(47) <= FROM_WINDOW_DEC_MASK(11);
UNWINDOWED_MASK(48) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(12);
UNWINDOWED_MASK(49) <= FROM_WINDOW_DEC_MASK(12);
UNWINDOWED_MASK(50) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(12);
UNWINDOWED_MASK(51) <= FROM_WINDOW_DEC_MASK(12);
UNWINDOWED_MASK(52) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(13);
UNWINDOWED_MASK(53) <= FROM_WINDOW_DEC_MASK(13);
UNWINDOWED_MASK(54) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(13);
UNWINDOWED_MASK(55) <= FROM_WINDOW_DEC_MASK(13);
UNWINDOWED_MASK(56) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(14);
UNWINDOWED_MASK(57) <= FROM_WINDOW_DEC_MASK(14);
UNWINDOWED_MASK(58) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(14);
UNWINDOWED_MASK(59) <= FROM_WINDOW_DEC_MASK(14);
UNWINDOWED_MASK(60) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(15);
UNWINDOWED_MASK(61) <= FROM_WINDOW_DEC_MASK(15);
UNWINDOWED_MASK(62) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(15);
UNWINDOWED_MASK(63) <= FROM_WINDOW_DEC_MASK(15);
UNWINDOWED_MASK(64) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(16);
UNWINDOWED_MASK(65) <= FROM_WINDOW_DEC_MASK(16);
UNWINDOWED_MASK(66) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(16);
UNWINDOWED_MASK(67) <= FROM_WINDOW_DEC_MASK(16);
UNWINDOWED_MASK(68) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(17);
UNWINDOWED_MASK(69) <= FROM_WINDOW_DEC_MASK(17);
UNWINDOWED_MASK(70) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(17);
UNWINDOWED_MASK(71) <= FROM_WINDOW_DEC_MASK(17);
UNWINDOWED_MASK(72) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(18);
UNWINDOWED_MASK(73) <= FROM_WINDOW_DEC_MASK(18);
UNWINDOWED_MASK(74) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(18);
UNWINDOWED_MASK(75) <= FROM_WINDOW_DEC_MASK(18);
UNWINDOWED_MASK(76) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(19);
UNWINDOWED_MASK(77) <= FROM_WINDOW_DEC_MASK(19);
UNWINDOWED_MASK(78) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(19);
UNWINDOWED_MASK(79) <= FROM_WINDOW_DEC_MASK(19);
UNWINDOWED_MASK(80) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(20);
UNWINDOWED_MASK(81) <= FROM_WINDOW_DEC_MASK(20);
UNWINDOWED_MASK(82) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(20);
UNWINDOWED_MASK(83) <= FROM_WINDOW_DEC_MASK(20);
UNWINDOWED_MASK(84) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(21);
UNWINDOWED_MASK(85) <= FROM_WINDOW_DEC_MASK(21);
UNWINDOWED_MASK(86) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(21);
UNWINDOWED_MASK(87) <= FROM_WINDOW_DEC_MASK(21);
UNWINDOWED_MASK(88) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(22);
UNWINDOWED_MASK(89) <= FROM_WINDOW_DEC_MASK(22);
UNWINDOWED_MASK(90) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(22);
UNWINDOWED_MASK(91) <= FROM_WINDOW_DEC_MASK(22);
UNWINDOWED_MASK(92) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(23);
UNWINDOWED_MASK(93) <= FROM_WINDOW_DEC_MASK(23);
UNWINDOWED_MASK(94) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(23);
UNWINDOWED_MASK(95) <= FROM_WINDOW_DEC_MASK(23);
UNWINDOWED_MASK(96) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(24);
UNWINDOWED_MASK(97) <= FROM_WINDOW_DEC_MASK(24);
UNWINDOWED_MASK(98) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(24);
UNWINDOWED_MASK(99) <= FROM_WINDOW_DEC_MASK(24);
UNWINDOWED_MASK(100) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(25);
UNWINDOWED_MASK(101) <= FROM_WINDOW_DEC_MASK(25);
UNWINDOWED_MASK(102) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(25);
UNWINDOWED_MASK(103) <= FROM_WINDOW_DEC_MASK(25);
UNWINDOWED_MASK(104) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(26);
UNWINDOWED_MASK(105) <= FROM_WINDOW_DEC_MASK(26);
UNWINDOWED_MASK(106) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(26);
UNWINDOWED_MASK(107) <= FROM_WINDOW_DEC_MASK(26);
UNWINDOWED_MASK(108) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(27);
UNWINDOWED_MASK(109) <= FROM_WINDOW_DEC_MASK(27);
UNWINDOWED_MASK(110) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(27);
UNWINDOWED_MASK(111) <= FROM_WINDOW_DEC_MASK(27);
UNWINDOWED_MASK(112) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(28);
UNWINDOWED_MASK(113) <= FROM_WINDOW_DEC_MASK(28);
UNWINDOWED_MASK(114) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(28);
UNWINDOWED_MASK(115) <= FROM_WINDOW_DEC_MASK(28);
UNWINDOWED_MASK(116) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(29);
UNWINDOWED_MASK(117) <= FROM_WINDOW_DEC_MASK(29);
UNWINDOWED_MASK(118) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(29);
UNWINDOWED_MASK(119) <= FROM_WINDOW_DEC_MASK(29);
UNWINDOWED_MASK(120) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(30);
UNWINDOWED_MASK(121) <= FROM_WINDOW_DEC_MASK(30);
UNWINDOWED_MASK(122) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(30);
UNWINDOWED_MASK(123) <= FROM_WINDOW_DEC_MASK(30);
UNWINDOWED_MASK(124) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(31);
UNWINDOWED_MASK(125) <= FROM_WINDOW_DEC_MASK(31);
UNWINDOWED_MASK(126) <= QEP_N_7_W_5_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(31);
UNWINDOWED_MASK(127) <= FROM_WINDOW_DEC_MASK(31);
UNWINDOWED_MASK(127) <= FROM_WINDOW_DEC_MASK(31);
MUX_REORD_UPDATE_0 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(0 DOWNTO 0) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(0 DOWNTO 0)
									);
MUX_REORD_UPDATE_1 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(2 DOWNTO 2) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(1 DOWNTO 1)
									);
MUX_REORD_UPDATE_2 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(4 DOWNTO 4) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(2 DOWNTO 2)
									);
MUX_REORD_UPDATE_3 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(6 DOWNTO 6) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(3 DOWNTO 3)
									);
MUX_REORD_UPDATE_4 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(8 DOWNTO 8) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(4 DOWNTO 4)
									);
MUX_REORD_UPDATE_5 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(10 DOWNTO 10) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(5 DOWNTO 5)
									);
MUX_REORD_UPDATE_6 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(12 DOWNTO 12) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(6 DOWNTO 6)
									);
MUX_REORD_UPDATE_7 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(14 DOWNTO 14) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(7 DOWNTO 7)
									);
MUX_REORD_UPDATE_8 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(16 DOWNTO 16) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(8 DOWNTO 8)
									);
MUX_REORD_UPDATE_9 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(18 DOWNTO 18) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(9 DOWNTO 9)
									);
MUX_REORD_UPDATE_10 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(20 DOWNTO 20) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(10 DOWNTO 10)
									);
MUX_REORD_UPDATE_11 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(22 DOWNTO 22) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(11 DOWNTO 11)
									);
MUX_REORD_UPDATE_12 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(24 DOWNTO 24) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(12 DOWNTO 12)
									);
MUX_REORD_UPDATE_13 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(26 DOWNTO 26) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(13 DOWNTO 13)
									);
MUX_REORD_UPDATE_14 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(28 DOWNTO 28) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(14 DOWNTO 14)
									);
MUX_REORD_UPDATE_15 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(30 DOWNTO 30) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(15 DOWNTO 15)
									);
MUX_REORD_UPDATE_16 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(32 DOWNTO 32) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(16 DOWNTO 16)
									);
MUX_REORD_UPDATE_17 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(34 DOWNTO 34) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(17 DOWNTO 17)
									);
MUX_REORD_UPDATE_18 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(36 DOWNTO 36) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(18 DOWNTO 18)
									);
MUX_REORD_UPDATE_19 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(38 DOWNTO 38) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(19 DOWNTO 19)
									);
MUX_REORD_UPDATE_20 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(40 DOWNTO 40) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(20 DOWNTO 20)
									);
MUX_REORD_UPDATE_21 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(42 DOWNTO 42) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(21 DOWNTO 21)
									);
MUX_REORD_UPDATE_22 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(44 DOWNTO 44) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(22 DOWNTO 22)
									);
MUX_REORD_UPDATE_23 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(46 DOWNTO 46) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(23 DOWNTO 23)
									);
MUX_REORD_UPDATE_24 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(48 DOWNTO 48) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(24 DOWNTO 24)
									);
MUX_REORD_UPDATE_25 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(50 DOWNTO 50) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(25 DOWNTO 25)
									);
MUX_REORD_UPDATE_26 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(52 DOWNTO 52) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(26 DOWNTO 26)
									);
MUX_REORD_UPDATE_27 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(54 DOWNTO 54) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(27 DOWNTO 27)
									);
MUX_REORD_UPDATE_28 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(56 DOWNTO 56) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(28 DOWNTO 28)
									);
MUX_REORD_UPDATE_29 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(58 DOWNTO 58) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(29 DOWNTO 29)
									);
MUX_REORD_UPDATE_30 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(60 DOWNTO 60) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(30 DOWNTO 30)
									);
MUX_REORD_UPDATE_31 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(62 DOWNTO 62) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(31 DOWNTO 31)
									);
MUX_REORD_UPDATE_32 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(64 DOWNTO 64) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(32 DOWNTO 32)
									);
MUX_REORD_UPDATE_33 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(66 DOWNTO 66) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(33 DOWNTO 33)
									);
MUX_REORD_UPDATE_34 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(68 DOWNTO 68) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(34 DOWNTO 34)
									);
MUX_REORD_UPDATE_35 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(70 DOWNTO 70) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(35 DOWNTO 35)
									);
MUX_REORD_UPDATE_36 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(72 DOWNTO 72) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(36 DOWNTO 36)
									);
MUX_REORD_UPDATE_37 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(74 DOWNTO 74) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(37 DOWNTO 37)
									);
MUX_REORD_UPDATE_38 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(76 DOWNTO 76) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(38 DOWNTO 38)
									);
MUX_REORD_UPDATE_39 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(78 DOWNTO 78) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(39 DOWNTO 39)
									);
MUX_REORD_UPDATE_40 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(80 DOWNTO 80) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(40 DOWNTO 40)
									);
MUX_REORD_UPDATE_41 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(82 DOWNTO 82) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(41 DOWNTO 41)
									);
MUX_REORD_UPDATE_42 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(84 DOWNTO 84) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(42 DOWNTO 42)
									);
MUX_REORD_UPDATE_43 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(86 DOWNTO 86) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(43 DOWNTO 43)
									);
MUX_REORD_UPDATE_44 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(88 DOWNTO 88) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(44 DOWNTO 44)
									);
MUX_REORD_UPDATE_45 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(90 DOWNTO 90) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(45 DOWNTO 45)
									);
MUX_REORD_UPDATE_46 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(92 DOWNTO 92) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(46 DOWNTO 46)
									);
MUX_REORD_UPDATE_47 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(94 DOWNTO 94) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(47 DOWNTO 47)
									);
MUX_REORD_UPDATE_48 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(96 DOWNTO 96) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(48 DOWNTO 48)
									);
MUX_REORD_UPDATE_49 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(98 DOWNTO 98) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(49 DOWNTO 49)
									);
MUX_REORD_UPDATE_50 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(100 DOWNTO 100) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(50 DOWNTO 50)
									);
MUX_REORD_UPDATE_51 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(102 DOWNTO 102) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(51 DOWNTO 51)
									);
MUX_REORD_UPDATE_52 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(104 DOWNTO 104) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(52 DOWNTO 52)
									);
MUX_REORD_UPDATE_53 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(106 DOWNTO 106) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(53 DOWNTO 53)
									);
MUX_REORD_UPDATE_54 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(108 DOWNTO 108) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(54 DOWNTO 54)
									);
MUX_REORD_UPDATE_55 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(110 DOWNTO 110) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(55 DOWNTO 55)
									);
MUX_REORD_UPDATE_56 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(112 DOWNTO 112) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(56 DOWNTO 56)
									);
MUX_REORD_UPDATE_57 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(114 DOWNTO 114) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(57 DOWNTO 57)
									);
MUX_REORD_UPDATE_58 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(116 DOWNTO 116) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(58 DOWNTO 58)
									);
MUX_REORD_UPDATE_59 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(118 DOWNTO 118) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(59 DOWNTO 59)
									);
MUX_REORD_UPDATE_60 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(120 DOWNTO 120) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(60 DOWNTO 60)
									);
MUX_REORD_UPDATE_61 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(122 DOWNTO 122) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(61 DOWNTO 61)
									);
MUX_REORD_UPDATE_62 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(124 DOWNTO 124) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(62 DOWNTO 62)
									);
MUX_REORD_UPDATE_63 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(126 DOWNTO 126) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(63 DOWNTO 63)
									);
MUX_REORD_UPDATE_64 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(64 DOWNTO 64) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(1 DOWNTO 1) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(64 DOWNTO 64)
									);
MUX_REORD_UPDATE_65 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(3 DOWNTO 3) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(65 DOWNTO 65)
									);
MUX_REORD_UPDATE_66 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(66 DOWNTO 66) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(5 DOWNTO 5) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(66 DOWNTO 66)
									);
MUX_REORD_UPDATE_67 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(7 DOWNTO 7) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(67 DOWNTO 67)
									);
MUX_REORD_UPDATE_68 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(68 DOWNTO 68) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(9 DOWNTO 9) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(68 DOWNTO 68)
									);
MUX_REORD_UPDATE_69 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(11 DOWNTO 11) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(69 DOWNTO 69)
									);
MUX_REORD_UPDATE_70 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(70 DOWNTO 70) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(13 DOWNTO 13) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(70 DOWNTO 70)
									);
MUX_REORD_UPDATE_71 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(15 DOWNTO 15) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(71 DOWNTO 71)
									);
MUX_REORD_UPDATE_72 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(72 DOWNTO 72) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(17 DOWNTO 17) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(72 DOWNTO 72)
									);
MUX_REORD_UPDATE_73 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(19 DOWNTO 19) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(73 DOWNTO 73)
									);
MUX_REORD_UPDATE_74 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(74 DOWNTO 74) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(21 DOWNTO 21) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(74 DOWNTO 74)
									);
MUX_REORD_UPDATE_75 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(23 DOWNTO 23) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(75 DOWNTO 75)
									);
MUX_REORD_UPDATE_76 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(76 DOWNTO 76) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(25 DOWNTO 25) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(76 DOWNTO 76)
									);
MUX_REORD_UPDATE_77 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(27 DOWNTO 27) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(77 DOWNTO 77)
									);
MUX_REORD_UPDATE_78 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(78 DOWNTO 78) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(29 DOWNTO 29) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(78 DOWNTO 78)
									);
MUX_REORD_UPDATE_79 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(31 DOWNTO 31) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(79 DOWNTO 79)
									);
MUX_REORD_UPDATE_80 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(80 DOWNTO 80) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(33 DOWNTO 33) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(80 DOWNTO 80)
									);
MUX_REORD_UPDATE_81 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(35 DOWNTO 35) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(81 DOWNTO 81)
									);
MUX_REORD_UPDATE_82 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(82 DOWNTO 82) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(37 DOWNTO 37) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(82 DOWNTO 82)
									);
MUX_REORD_UPDATE_83 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(39 DOWNTO 39) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(83 DOWNTO 83)
									);
MUX_REORD_UPDATE_84 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(84 DOWNTO 84) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(41 DOWNTO 41) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(84 DOWNTO 84)
									);
MUX_REORD_UPDATE_85 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(43 DOWNTO 43) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(85 DOWNTO 85)
									);
MUX_REORD_UPDATE_86 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(86 DOWNTO 86) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(45 DOWNTO 45) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(86 DOWNTO 86)
									);
MUX_REORD_UPDATE_87 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(47 DOWNTO 47) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(87 DOWNTO 87)
									);
MUX_REORD_UPDATE_88 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(88 DOWNTO 88) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(49 DOWNTO 49) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(88 DOWNTO 88)
									);
MUX_REORD_UPDATE_89 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(51 DOWNTO 51) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(89 DOWNTO 89)
									);
MUX_REORD_UPDATE_90 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(90 DOWNTO 90) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(53 DOWNTO 53) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(90 DOWNTO 90)
									);
MUX_REORD_UPDATE_91 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(55 DOWNTO 55) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(91 DOWNTO 91)
									);
MUX_REORD_UPDATE_92 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(92 DOWNTO 92) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(57 DOWNTO 57) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(92 DOWNTO 92)
									);
MUX_REORD_UPDATE_93 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(59 DOWNTO 59) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(93 DOWNTO 93)
									);
MUX_REORD_UPDATE_94 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(94 DOWNTO 94) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(61 DOWNTO 61) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(94 DOWNTO 94)
									);
MUX_REORD_UPDATE_95 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(63 DOWNTO 63) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(95 DOWNTO 95)
									);
MUX_REORD_UPDATE_96 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(96 DOWNTO 96) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(65 DOWNTO 65) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(65 DOWNTO 65) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(96 DOWNTO 96)
									);
MUX_REORD_UPDATE_97 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(67 DOWNTO 67) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(67 DOWNTO 67) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(97 DOWNTO 97)
									);
MUX_REORD_UPDATE_98 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(98 DOWNTO 98) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(69 DOWNTO 69) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(69 DOWNTO 69) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(98 DOWNTO 98)
									);
MUX_REORD_UPDATE_99 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(71 DOWNTO 71) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(71 DOWNTO 71) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(99 DOWNTO 99)
									);
MUX_REORD_UPDATE_100 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(100 DOWNTO 100) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(73 DOWNTO 73) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(73 DOWNTO 73) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(100 DOWNTO 100)
									);
MUX_REORD_UPDATE_101 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(75 DOWNTO 75) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(75 DOWNTO 75) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(101 DOWNTO 101)
									);
MUX_REORD_UPDATE_102 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(102 DOWNTO 102) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(77 DOWNTO 77) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(77 DOWNTO 77) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(102 DOWNTO 102)
									);
MUX_REORD_UPDATE_103 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(79 DOWNTO 79) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(79 DOWNTO 79) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(103 DOWNTO 103)
									);
MUX_REORD_UPDATE_104 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(104 DOWNTO 104) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(81 DOWNTO 81) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(81 DOWNTO 81) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(104 DOWNTO 104)
									);
MUX_REORD_UPDATE_105 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(83 DOWNTO 83) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(83 DOWNTO 83) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(105 DOWNTO 105)
									);
MUX_REORD_UPDATE_106 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(106 DOWNTO 106) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(85 DOWNTO 85) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(85 DOWNTO 85) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(106 DOWNTO 106)
									);
MUX_REORD_UPDATE_107 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(87 DOWNTO 87) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(87 DOWNTO 87) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(107 DOWNTO 107)
									);
MUX_REORD_UPDATE_108 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(108 DOWNTO 108) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(89 DOWNTO 89) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(89 DOWNTO 89) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(108 DOWNTO 108)
									);
MUX_REORD_UPDATE_109 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(91 DOWNTO 91) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(91 DOWNTO 91) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(109 DOWNTO 109)
									);
MUX_REORD_UPDATE_110 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(110 DOWNTO 110) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(93 DOWNTO 93) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(93 DOWNTO 93) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(110 DOWNTO 110)
									);
MUX_REORD_UPDATE_111 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(95 DOWNTO 95) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(95 DOWNTO 95) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(111 DOWNTO 111)
									);
MUX_REORD_UPDATE_112 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(112 DOWNTO 112) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(97 DOWNTO 97) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(97 DOWNTO 97) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(112 DOWNTO 112)
									);
MUX_REORD_UPDATE_113 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(99 DOWNTO 99) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(99 DOWNTO 99) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(113 DOWNTO 113)
									);
MUX_REORD_UPDATE_114 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(114 DOWNTO 114) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(101 DOWNTO 101) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(101 DOWNTO 101) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(114 DOWNTO 114)
									);
MUX_REORD_UPDATE_115 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(103 DOWNTO 103) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(103 DOWNTO 103) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(115 DOWNTO 115)
									);
MUX_REORD_UPDATE_116 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(116 DOWNTO 116) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(105 DOWNTO 105) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(105 DOWNTO 105) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(116 DOWNTO 116)
									);
MUX_REORD_UPDATE_117 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(107 DOWNTO 107) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(107 DOWNTO 107) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(117 DOWNTO 117)
									);
MUX_REORD_UPDATE_118 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(118 DOWNTO 118) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(109 DOWNTO 109) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(109 DOWNTO 109) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(118 DOWNTO 118)
									);
MUX_REORD_UPDATE_119 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(111 DOWNTO 111) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(111 DOWNTO 111) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(119 DOWNTO 119)
									);
MUX_REORD_UPDATE_120 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(120 DOWNTO 120) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(113 DOWNTO 113) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(113 DOWNTO 113) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(120 DOWNTO 120)
									);
MUX_REORD_UPDATE_121 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(115 DOWNTO 115) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(115 DOWNTO 115) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(121 DOWNTO 121)
									);
MUX_REORD_UPDATE_122 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(122 DOWNTO 122) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(117 DOWNTO 117) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(117 DOWNTO 117) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(122 DOWNTO 122)
									);
MUX_REORD_UPDATE_123 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(119 DOWNTO 119) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(119 DOWNTO 119) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(123 DOWNTO 123)
									);
MUX_REORD_UPDATE_124 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(124 DOWNTO 124) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(121 DOWNTO 121) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(121 DOWNTO 121) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(124 DOWNTO 124)
									);
MUX_REORD_UPDATE_125 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(123 DOWNTO 123) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(123 DOWNTO 123) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(125 DOWNTO 125)
									);
MUX_REORD_UPDATE_126 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(126 DOWNTO 126) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(125 DOWNTO 125) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(125 DOWNTO 125) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(126 DOWNTO 126)
									);
MUX_REORD_UPDATE_127 : multiplexer_7_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_7_1_IN_1 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_7_1_IN_2 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_7_1_IN_3 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_7_1_IN_4 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_7_1_IN_5 => UNWINDOWED_MASK(127 DOWNTO 127) ,
										MUX_7_1_IN_6 => UNWINDOWED_MASK(127 DOWNTO 127) ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => REORDERED_MASK(127 DOWNTO 127)
									);

STATE_UPDATE_MASK(0) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(0) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(0);
STATE_UPDATE_MASK(1) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(1);
STATE_UPDATE_MASK(2) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(2) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(2);
STATE_UPDATE_MASK(3) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(3) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(3);
STATE_UPDATE_MASK(4) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(4) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(4);
STATE_UPDATE_MASK(5) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(5) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(5);
STATE_UPDATE_MASK(6) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(6) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(6);
STATE_UPDATE_MASK(7) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(7) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(7);
STATE_UPDATE_MASK(8) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(8) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(8);
STATE_UPDATE_MASK(9) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(9) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(9);
STATE_UPDATE_MASK(10) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(10) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(10);
STATE_UPDATE_MASK(11) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(11) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(11);
STATE_UPDATE_MASK(12) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(12) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(12);
STATE_UPDATE_MASK(13) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(13) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(13);
STATE_UPDATE_MASK(14) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(14) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(14);
STATE_UPDATE_MASK(15) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(15) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(15);
STATE_UPDATE_MASK(16) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(16) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(16);
STATE_UPDATE_MASK(17) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(17) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(17);
STATE_UPDATE_MASK(18) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(18) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(18);
STATE_UPDATE_MASK(19) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(19) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(19);
STATE_UPDATE_MASK(20) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(20) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(20);
STATE_UPDATE_MASK(21) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(21) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(21);
STATE_UPDATE_MASK(22) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(22) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(22);
STATE_UPDATE_MASK(23) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(23) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(23);
STATE_UPDATE_MASK(24) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(24) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(24);
STATE_UPDATE_MASK(25) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(25) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(25);
STATE_UPDATE_MASK(26) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(26) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(26);
STATE_UPDATE_MASK(27) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(27) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(27);
STATE_UPDATE_MASK(28) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(28) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(28);
STATE_UPDATE_MASK(29) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(29) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(29);
STATE_UPDATE_MASK(30) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(30) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(30);
STATE_UPDATE_MASK(31) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(31) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(31);
STATE_UPDATE_MASK(32) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(32) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(32);
STATE_UPDATE_MASK(33) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(33) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(33);
STATE_UPDATE_MASK(34) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(34) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(34);
STATE_UPDATE_MASK(35) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(35) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(35);
STATE_UPDATE_MASK(36) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(36) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(36);
STATE_UPDATE_MASK(37) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(37) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(37);
STATE_UPDATE_MASK(38) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(38) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(38);
STATE_UPDATE_MASK(39) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(39) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(39);
STATE_UPDATE_MASK(40) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(40) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(40);
STATE_UPDATE_MASK(41) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(41) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(41);
STATE_UPDATE_MASK(42) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(42) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(42);
STATE_UPDATE_MASK(43) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(43) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(43);
STATE_UPDATE_MASK(44) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(44) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(44);
STATE_UPDATE_MASK(45) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(45) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(45);
STATE_UPDATE_MASK(46) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(46) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(46);
STATE_UPDATE_MASK(47) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(47) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(47);
STATE_UPDATE_MASK(48) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(48) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(48);
STATE_UPDATE_MASK(49) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(49) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(49);
STATE_UPDATE_MASK(50) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(50) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(50);
STATE_UPDATE_MASK(51) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(51) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(51);
STATE_UPDATE_MASK(52) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(52) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(52);
STATE_UPDATE_MASK(53) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(53) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(53);
STATE_UPDATE_MASK(54) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(54) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(54);
STATE_UPDATE_MASK(55) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(55) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(55);
STATE_UPDATE_MASK(56) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(56) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(56);
STATE_UPDATE_MASK(57) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(57) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(57);
STATE_UPDATE_MASK(58) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(58) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(58);
STATE_UPDATE_MASK(59) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(59) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(59);
STATE_UPDATE_MASK(60) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(60) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(60);
STATE_UPDATE_MASK(61) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(61) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(61);
STATE_UPDATE_MASK(62) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(62) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(62);
STATE_UPDATE_MASK(63) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(63) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(63);
STATE_UPDATE_MASK(64) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(64) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(64);
STATE_UPDATE_MASK(65) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(65) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(65);
STATE_UPDATE_MASK(66) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(66) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(66);
STATE_UPDATE_MASK(67) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(67) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(67);
STATE_UPDATE_MASK(68) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(68) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(68);
STATE_UPDATE_MASK(69) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(69) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(69);
STATE_UPDATE_MASK(70) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(70) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(70);
STATE_UPDATE_MASK(71) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(71) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(71);
STATE_UPDATE_MASK(72) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(72) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(72);
STATE_UPDATE_MASK(73) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(73) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(73);
STATE_UPDATE_MASK(74) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(74) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(74);
STATE_UPDATE_MASK(75) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(75) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(75);
STATE_UPDATE_MASK(76) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(76) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(76);
STATE_UPDATE_MASK(77) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(77) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(77);
STATE_UPDATE_MASK(78) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(78) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(78);
STATE_UPDATE_MASK(79) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(79) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(79);
STATE_UPDATE_MASK(80) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(80) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(80);
STATE_UPDATE_MASK(81) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(81) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(81);
STATE_UPDATE_MASK(82) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(82) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(82);
STATE_UPDATE_MASK(83) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(83) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(83);
STATE_UPDATE_MASK(84) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(84) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(84);
STATE_UPDATE_MASK(85) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(85) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(85);
STATE_UPDATE_MASK(86) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(86) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(86);
STATE_UPDATE_MASK(87) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(87) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(87);
STATE_UPDATE_MASK(88) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(88) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(88);
STATE_UPDATE_MASK(89) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(89) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(89);
STATE_UPDATE_MASK(90) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(90) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(90);
STATE_UPDATE_MASK(91) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(91) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(91);
STATE_UPDATE_MASK(92) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(92) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(92);
STATE_UPDATE_MASK(93) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(93) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(93);
STATE_UPDATE_MASK(94) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(94) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(94);
STATE_UPDATE_MASK(95) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(95) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(95);
STATE_UPDATE_MASK(96) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(96) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(96);
STATE_UPDATE_MASK(97) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(97) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(97);
STATE_UPDATE_MASK(98) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(98) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(98);
STATE_UPDATE_MASK(99) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(99) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(99);
STATE_UPDATE_MASK(100) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(100) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(100);
STATE_UPDATE_MASK(101) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(101) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(101);
STATE_UPDATE_MASK(102) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(102) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(102);
STATE_UPDATE_MASK(103) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(103) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(103);
STATE_UPDATE_MASK(104) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(104) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(104);
STATE_UPDATE_MASK(105) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(105) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(105);
STATE_UPDATE_MASK(106) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(106) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(106);
STATE_UPDATE_MASK(107) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(107) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(107);
STATE_UPDATE_MASK(108) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(108) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(108);
STATE_UPDATE_MASK(109) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(109) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(109);
STATE_UPDATE_MASK(110) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(110) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(110);
STATE_UPDATE_MASK(111) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(111) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(111);
STATE_UPDATE_MASK(112) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(112) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(112);
STATE_UPDATE_MASK(113) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(113) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(113);
STATE_UPDATE_MASK(114) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(114) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(114);
STATE_UPDATE_MASK(115) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(115) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(115);
STATE_UPDATE_MASK(116) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(116) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(116);
STATE_UPDATE_MASK(117) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(117) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(117);
STATE_UPDATE_MASK(118) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(118) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(118);
STATE_UPDATE_MASK(119) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(119) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(119);
STATE_UPDATE_MASK(120) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(120) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(120);
STATE_UPDATE_MASK(121) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(121) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(121);
STATE_UPDATE_MASK(122) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(122) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(122);
STATE_UPDATE_MASK(123) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(123) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(123);
STATE_UPDATE_MASK(124) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(124) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(124);
STATE_UPDATE_MASK(125) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(125) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(125);
STATE_UPDATE_MASK(126) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(126) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(126);
STATE_UPDATE_MASK(127) <= QEP_N_7_W_5_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(127) AND QEP_N_7_W_5_S_0_IN_CTRL_MASK(127);

QEP_N_7_W_5_S_0_OUT_DONE <= FROM_FIRST_CU_DONE;
CONTROL_UNIT_0 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_7_W_5_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_7_W_5_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
		CONTROL_UNIT_OUT_DONE => FROM_FIRST_CU_DONE );
CONTROL_UNIT_1 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_7_W_5_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_7_W_5_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0));

DATAPATH_0: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_0 ,
            DATAPATH_IN_B => FROM_WINDOW_1 ,
            DATAPATH_IN_SINE => QEP_N_7_W_5_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_7_W_5_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_0 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1);
DATAPATH_1: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_2 ,
            DATAPATH_IN_B => FROM_WINDOW_3 ,
            DATAPATH_IN_SINE => QEP_N_7_W_5_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_7_W_5_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_7_W_5_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_7_W_5_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_2 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_3);

UNWINDOWED_0 <= FROM_DATAPATHS_0;
UNWINDOWED_1 <= FROM_DATAPATHS_1;
UNWINDOWED_2 <= FROM_DATAPATHS_2;
UNWINDOWED_3 <= FROM_DATAPATHS_3;
UNWINDOWED_4 <= FROM_DATAPATHS_0;
UNWINDOWED_5 <= FROM_DATAPATHS_1;
UNWINDOWED_6 <= FROM_DATAPATHS_2;
UNWINDOWED_7 <= FROM_DATAPATHS_3;
UNWINDOWED_8 <= FROM_DATAPATHS_0;
UNWINDOWED_9 <= FROM_DATAPATHS_1;
UNWINDOWED_10 <= FROM_DATAPATHS_2;
UNWINDOWED_11 <= FROM_DATAPATHS_3;
UNWINDOWED_12 <= FROM_DATAPATHS_0;
UNWINDOWED_13 <= FROM_DATAPATHS_1;
UNWINDOWED_14 <= FROM_DATAPATHS_2;
UNWINDOWED_15 <= FROM_DATAPATHS_3;
UNWINDOWED_16 <= FROM_DATAPATHS_0;
UNWINDOWED_17 <= FROM_DATAPATHS_1;
UNWINDOWED_18 <= FROM_DATAPATHS_2;
UNWINDOWED_19 <= FROM_DATAPATHS_3;
UNWINDOWED_20 <= FROM_DATAPATHS_0;
UNWINDOWED_21 <= FROM_DATAPATHS_1;
UNWINDOWED_22 <= FROM_DATAPATHS_2;
UNWINDOWED_23 <= FROM_DATAPATHS_3;
UNWINDOWED_24 <= FROM_DATAPATHS_0;
UNWINDOWED_25 <= FROM_DATAPATHS_1;
UNWINDOWED_26 <= FROM_DATAPATHS_2;
UNWINDOWED_27 <= FROM_DATAPATHS_3;
UNWINDOWED_28 <= FROM_DATAPATHS_0;
UNWINDOWED_29 <= FROM_DATAPATHS_1;
UNWINDOWED_30 <= FROM_DATAPATHS_2;
UNWINDOWED_31 <= FROM_DATAPATHS_3;
UNWINDOWED_32 <= FROM_DATAPATHS_0;
UNWINDOWED_33 <= FROM_DATAPATHS_1;
UNWINDOWED_34 <= FROM_DATAPATHS_2;
UNWINDOWED_35 <= FROM_DATAPATHS_3;
UNWINDOWED_36 <= FROM_DATAPATHS_0;
UNWINDOWED_37 <= FROM_DATAPATHS_1;
UNWINDOWED_38 <= FROM_DATAPATHS_2;
UNWINDOWED_39 <= FROM_DATAPATHS_3;
UNWINDOWED_40 <= FROM_DATAPATHS_0;
UNWINDOWED_41 <= FROM_DATAPATHS_1;
UNWINDOWED_42 <= FROM_DATAPATHS_2;
UNWINDOWED_43 <= FROM_DATAPATHS_3;
UNWINDOWED_44 <= FROM_DATAPATHS_0;
UNWINDOWED_45 <= FROM_DATAPATHS_1;
UNWINDOWED_46 <= FROM_DATAPATHS_2;
UNWINDOWED_47 <= FROM_DATAPATHS_3;
UNWINDOWED_48 <= FROM_DATAPATHS_0;
UNWINDOWED_49 <= FROM_DATAPATHS_1;
UNWINDOWED_50 <= FROM_DATAPATHS_2;
UNWINDOWED_51 <= FROM_DATAPATHS_3;
UNWINDOWED_52 <= FROM_DATAPATHS_0;
UNWINDOWED_53 <= FROM_DATAPATHS_1;
UNWINDOWED_54 <= FROM_DATAPATHS_2;
UNWINDOWED_55 <= FROM_DATAPATHS_3;
UNWINDOWED_56 <= FROM_DATAPATHS_0;
UNWINDOWED_57 <= FROM_DATAPATHS_1;
UNWINDOWED_58 <= FROM_DATAPATHS_2;
UNWINDOWED_59 <= FROM_DATAPATHS_3;
UNWINDOWED_60 <= FROM_DATAPATHS_0;
UNWINDOWED_61 <= FROM_DATAPATHS_1;
UNWINDOWED_62 <= FROM_DATAPATHS_2;
UNWINDOWED_63 <= FROM_DATAPATHS_3;
UNWINDOWED_64 <= FROM_DATAPATHS_0;
UNWINDOWED_65 <= FROM_DATAPATHS_1;
UNWINDOWED_66 <= FROM_DATAPATHS_2;
UNWINDOWED_67 <= FROM_DATAPATHS_3;
UNWINDOWED_68 <= FROM_DATAPATHS_0;
UNWINDOWED_69 <= FROM_DATAPATHS_1;
UNWINDOWED_70 <= FROM_DATAPATHS_2;
UNWINDOWED_71 <= FROM_DATAPATHS_3;
UNWINDOWED_72 <= FROM_DATAPATHS_0;
UNWINDOWED_73 <= FROM_DATAPATHS_1;
UNWINDOWED_74 <= FROM_DATAPATHS_2;
UNWINDOWED_75 <= FROM_DATAPATHS_3;
UNWINDOWED_76 <= FROM_DATAPATHS_0;
UNWINDOWED_77 <= FROM_DATAPATHS_1;
UNWINDOWED_78 <= FROM_DATAPATHS_2;
UNWINDOWED_79 <= FROM_DATAPATHS_3;
UNWINDOWED_80 <= FROM_DATAPATHS_0;
UNWINDOWED_81 <= FROM_DATAPATHS_1;
UNWINDOWED_82 <= FROM_DATAPATHS_2;
UNWINDOWED_83 <= FROM_DATAPATHS_3;
UNWINDOWED_84 <= FROM_DATAPATHS_0;
UNWINDOWED_85 <= FROM_DATAPATHS_1;
UNWINDOWED_86 <= FROM_DATAPATHS_2;
UNWINDOWED_87 <= FROM_DATAPATHS_3;
UNWINDOWED_88 <= FROM_DATAPATHS_0;
UNWINDOWED_89 <= FROM_DATAPATHS_1;
UNWINDOWED_90 <= FROM_DATAPATHS_2;
UNWINDOWED_91 <= FROM_DATAPATHS_3;
UNWINDOWED_92 <= FROM_DATAPATHS_0;
UNWINDOWED_93 <= FROM_DATAPATHS_1;
UNWINDOWED_94 <= FROM_DATAPATHS_2;
UNWINDOWED_95 <= FROM_DATAPATHS_3;
UNWINDOWED_96 <= FROM_DATAPATHS_0;
UNWINDOWED_97 <= FROM_DATAPATHS_1;
UNWINDOWED_98 <= FROM_DATAPATHS_2;
UNWINDOWED_99 <= FROM_DATAPATHS_3;
UNWINDOWED_100 <= FROM_DATAPATHS_0;
UNWINDOWED_101 <= FROM_DATAPATHS_1;
UNWINDOWED_102 <= FROM_DATAPATHS_2;
UNWINDOWED_103 <= FROM_DATAPATHS_3;
UNWINDOWED_104 <= FROM_DATAPATHS_0;
UNWINDOWED_105 <= FROM_DATAPATHS_1;
UNWINDOWED_106 <= FROM_DATAPATHS_2;
UNWINDOWED_107 <= FROM_DATAPATHS_3;
UNWINDOWED_108 <= FROM_DATAPATHS_0;
UNWINDOWED_109 <= FROM_DATAPATHS_1;
UNWINDOWED_110 <= FROM_DATAPATHS_2;
UNWINDOWED_111 <= FROM_DATAPATHS_3;
UNWINDOWED_112 <= FROM_DATAPATHS_0;
UNWINDOWED_113 <= FROM_DATAPATHS_1;
UNWINDOWED_114 <= FROM_DATAPATHS_2;
UNWINDOWED_115 <= FROM_DATAPATHS_3;
UNWINDOWED_116 <= FROM_DATAPATHS_0;
UNWINDOWED_117 <= FROM_DATAPATHS_1;
UNWINDOWED_118 <= FROM_DATAPATHS_2;
UNWINDOWED_119 <= FROM_DATAPATHS_3;
UNWINDOWED_120 <= FROM_DATAPATHS_0;
UNWINDOWED_121 <= FROM_DATAPATHS_1;
UNWINDOWED_122 <= FROM_DATAPATHS_2;
UNWINDOWED_123 <= FROM_DATAPATHS_3;
UNWINDOWED_124 <= FROM_DATAPATHS_0;
UNWINDOWED_125 <= FROM_DATAPATHS_1;
UNWINDOWED_126 <= FROM_DATAPATHS_2;
UNWINDOWED_127 <= FROM_DATAPATHS_3;

MUX_REORD_UNIT_0 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_0 ,
										MUX_7_1_IN_1 => UNWINDOWED_0 ,
										MUX_7_1_IN_2 => UNWINDOWED_0 ,
										MUX_7_1_IN_3 => UNWINDOWED_0 ,
										MUX_7_1_IN_4 => UNWINDOWED_0 ,
										MUX_7_1_IN_5 => UNWINDOWED_0 ,
										MUX_7_1_IN_6 => UNWINDOWED_0 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_0
									);
MUX_REORD_UNIT_1 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_1 ,
										MUX_7_1_IN_1 => UNWINDOWED_2 ,
										MUX_7_1_IN_2 => UNWINDOWED_2 ,
										MUX_7_1_IN_3 => UNWINDOWED_2 ,
										MUX_7_1_IN_4 => UNWINDOWED_2 ,
										MUX_7_1_IN_5 => UNWINDOWED_2 ,
										MUX_7_1_IN_6 => UNWINDOWED_2 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_1
									);
MUX_REORD_UNIT_2 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_2 ,
										MUX_7_1_IN_1 => UNWINDOWED_1 ,
										MUX_7_1_IN_2 => UNWINDOWED_4 ,
										MUX_7_1_IN_3 => UNWINDOWED_4 ,
										MUX_7_1_IN_4 => UNWINDOWED_4 ,
										MUX_7_1_IN_5 => UNWINDOWED_4 ,
										MUX_7_1_IN_6 => UNWINDOWED_4 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_2
									);
MUX_REORD_UNIT_3 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_3 ,
										MUX_7_1_IN_1 => UNWINDOWED_3 ,
										MUX_7_1_IN_2 => UNWINDOWED_6 ,
										MUX_7_1_IN_3 => UNWINDOWED_6 ,
										MUX_7_1_IN_4 => UNWINDOWED_6 ,
										MUX_7_1_IN_5 => UNWINDOWED_6 ,
										MUX_7_1_IN_6 => UNWINDOWED_6 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_3
									);
MUX_REORD_UNIT_4 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_4 ,
										MUX_7_1_IN_1 => UNWINDOWED_4 ,
										MUX_7_1_IN_2 => UNWINDOWED_1 ,
										MUX_7_1_IN_3 => UNWINDOWED_8 ,
										MUX_7_1_IN_4 => UNWINDOWED_8 ,
										MUX_7_1_IN_5 => UNWINDOWED_8 ,
										MUX_7_1_IN_6 => UNWINDOWED_8 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_4
									);
MUX_REORD_UNIT_5 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_5 ,
										MUX_7_1_IN_1 => UNWINDOWED_6 ,
										MUX_7_1_IN_2 => UNWINDOWED_3 ,
										MUX_7_1_IN_3 => UNWINDOWED_10 ,
										MUX_7_1_IN_4 => UNWINDOWED_10 ,
										MUX_7_1_IN_5 => UNWINDOWED_10 ,
										MUX_7_1_IN_6 => UNWINDOWED_10 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_5
									);
MUX_REORD_UNIT_6 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_6 ,
										MUX_7_1_IN_1 => UNWINDOWED_5 ,
										MUX_7_1_IN_2 => UNWINDOWED_5 ,
										MUX_7_1_IN_3 => UNWINDOWED_12 ,
										MUX_7_1_IN_4 => UNWINDOWED_12 ,
										MUX_7_1_IN_5 => UNWINDOWED_12 ,
										MUX_7_1_IN_6 => UNWINDOWED_12 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_6
									);
MUX_REORD_UNIT_7 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_7 ,
										MUX_7_1_IN_1 => UNWINDOWED_7 ,
										MUX_7_1_IN_2 => UNWINDOWED_7 ,
										MUX_7_1_IN_3 => UNWINDOWED_14 ,
										MUX_7_1_IN_4 => UNWINDOWED_14 ,
										MUX_7_1_IN_5 => UNWINDOWED_14 ,
										MUX_7_1_IN_6 => UNWINDOWED_14 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_7
									);
MUX_REORD_UNIT_8 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_8 ,
										MUX_7_1_IN_1 => UNWINDOWED_8 ,
										MUX_7_1_IN_2 => UNWINDOWED_8 ,
										MUX_7_1_IN_3 => UNWINDOWED_1 ,
										MUX_7_1_IN_4 => UNWINDOWED_16 ,
										MUX_7_1_IN_5 => UNWINDOWED_16 ,
										MUX_7_1_IN_6 => UNWINDOWED_16 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_8
									);
MUX_REORD_UNIT_9 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_9 ,
										MUX_7_1_IN_1 => UNWINDOWED_10 ,
										MUX_7_1_IN_2 => UNWINDOWED_10 ,
										MUX_7_1_IN_3 => UNWINDOWED_3 ,
										MUX_7_1_IN_4 => UNWINDOWED_18 ,
										MUX_7_1_IN_5 => UNWINDOWED_18 ,
										MUX_7_1_IN_6 => UNWINDOWED_18 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_9
									);
MUX_REORD_UNIT_10 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_10 ,
										MUX_7_1_IN_1 => UNWINDOWED_9 ,
										MUX_7_1_IN_2 => UNWINDOWED_12 ,
										MUX_7_1_IN_3 => UNWINDOWED_5 ,
										MUX_7_1_IN_4 => UNWINDOWED_20 ,
										MUX_7_1_IN_5 => UNWINDOWED_20 ,
										MUX_7_1_IN_6 => UNWINDOWED_20 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_10
									);
MUX_REORD_UNIT_11 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_11 ,
										MUX_7_1_IN_1 => UNWINDOWED_11 ,
										MUX_7_1_IN_2 => UNWINDOWED_14 ,
										MUX_7_1_IN_3 => UNWINDOWED_7 ,
										MUX_7_1_IN_4 => UNWINDOWED_22 ,
										MUX_7_1_IN_5 => UNWINDOWED_22 ,
										MUX_7_1_IN_6 => UNWINDOWED_22 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_11
									);
MUX_REORD_UNIT_12 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_12 ,
										MUX_7_1_IN_1 => UNWINDOWED_12 ,
										MUX_7_1_IN_2 => UNWINDOWED_9 ,
										MUX_7_1_IN_3 => UNWINDOWED_9 ,
										MUX_7_1_IN_4 => UNWINDOWED_24 ,
										MUX_7_1_IN_5 => UNWINDOWED_24 ,
										MUX_7_1_IN_6 => UNWINDOWED_24 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_12
									);
MUX_REORD_UNIT_13 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_13 ,
										MUX_7_1_IN_1 => UNWINDOWED_14 ,
										MUX_7_1_IN_2 => UNWINDOWED_11 ,
										MUX_7_1_IN_3 => UNWINDOWED_11 ,
										MUX_7_1_IN_4 => UNWINDOWED_26 ,
										MUX_7_1_IN_5 => UNWINDOWED_26 ,
										MUX_7_1_IN_6 => UNWINDOWED_26 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_13
									);
MUX_REORD_UNIT_14 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_14 ,
										MUX_7_1_IN_1 => UNWINDOWED_13 ,
										MUX_7_1_IN_2 => UNWINDOWED_13 ,
										MUX_7_1_IN_3 => UNWINDOWED_13 ,
										MUX_7_1_IN_4 => UNWINDOWED_28 ,
										MUX_7_1_IN_5 => UNWINDOWED_28 ,
										MUX_7_1_IN_6 => UNWINDOWED_28 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_14
									);
MUX_REORD_UNIT_15 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_15 ,
										MUX_7_1_IN_1 => UNWINDOWED_15 ,
										MUX_7_1_IN_2 => UNWINDOWED_15 ,
										MUX_7_1_IN_3 => UNWINDOWED_15 ,
										MUX_7_1_IN_4 => UNWINDOWED_30 ,
										MUX_7_1_IN_5 => UNWINDOWED_30 ,
										MUX_7_1_IN_6 => UNWINDOWED_30 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_15
									);
MUX_REORD_UNIT_16 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_16 ,
										MUX_7_1_IN_1 => UNWINDOWED_16 ,
										MUX_7_1_IN_2 => UNWINDOWED_16 ,
										MUX_7_1_IN_3 => UNWINDOWED_16 ,
										MUX_7_1_IN_4 => UNWINDOWED_1 ,
										MUX_7_1_IN_5 => UNWINDOWED_32 ,
										MUX_7_1_IN_6 => UNWINDOWED_32 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_16
									);
MUX_REORD_UNIT_17 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_17 ,
										MUX_7_1_IN_1 => UNWINDOWED_18 ,
										MUX_7_1_IN_2 => UNWINDOWED_18 ,
										MUX_7_1_IN_3 => UNWINDOWED_18 ,
										MUX_7_1_IN_4 => UNWINDOWED_3 ,
										MUX_7_1_IN_5 => UNWINDOWED_34 ,
										MUX_7_1_IN_6 => UNWINDOWED_34 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_17
									);
MUX_REORD_UNIT_18 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_18 ,
										MUX_7_1_IN_1 => UNWINDOWED_17 ,
										MUX_7_1_IN_2 => UNWINDOWED_20 ,
										MUX_7_1_IN_3 => UNWINDOWED_20 ,
										MUX_7_1_IN_4 => UNWINDOWED_5 ,
										MUX_7_1_IN_5 => UNWINDOWED_36 ,
										MUX_7_1_IN_6 => UNWINDOWED_36 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_18
									);
MUX_REORD_UNIT_19 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_19 ,
										MUX_7_1_IN_1 => UNWINDOWED_19 ,
										MUX_7_1_IN_2 => UNWINDOWED_22 ,
										MUX_7_1_IN_3 => UNWINDOWED_22 ,
										MUX_7_1_IN_4 => UNWINDOWED_7 ,
										MUX_7_1_IN_5 => UNWINDOWED_38 ,
										MUX_7_1_IN_6 => UNWINDOWED_38 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_19
									);
MUX_REORD_UNIT_20 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_20 ,
										MUX_7_1_IN_1 => UNWINDOWED_20 ,
										MUX_7_1_IN_2 => UNWINDOWED_17 ,
										MUX_7_1_IN_3 => UNWINDOWED_24 ,
										MUX_7_1_IN_4 => UNWINDOWED_9 ,
										MUX_7_1_IN_5 => UNWINDOWED_40 ,
										MUX_7_1_IN_6 => UNWINDOWED_40 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_20
									);
MUX_REORD_UNIT_21 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_21 ,
										MUX_7_1_IN_1 => UNWINDOWED_22 ,
										MUX_7_1_IN_2 => UNWINDOWED_19 ,
										MUX_7_1_IN_3 => UNWINDOWED_26 ,
										MUX_7_1_IN_4 => UNWINDOWED_11 ,
										MUX_7_1_IN_5 => UNWINDOWED_42 ,
										MUX_7_1_IN_6 => UNWINDOWED_42 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_21
									);
MUX_REORD_UNIT_22 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_22 ,
										MUX_7_1_IN_1 => UNWINDOWED_21 ,
										MUX_7_1_IN_2 => UNWINDOWED_21 ,
										MUX_7_1_IN_3 => UNWINDOWED_28 ,
										MUX_7_1_IN_4 => UNWINDOWED_13 ,
										MUX_7_1_IN_5 => UNWINDOWED_44 ,
										MUX_7_1_IN_6 => UNWINDOWED_44 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_22
									);
MUX_REORD_UNIT_23 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_23 ,
										MUX_7_1_IN_1 => UNWINDOWED_23 ,
										MUX_7_1_IN_2 => UNWINDOWED_23 ,
										MUX_7_1_IN_3 => UNWINDOWED_30 ,
										MUX_7_1_IN_4 => UNWINDOWED_15 ,
										MUX_7_1_IN_5 => UNWINDOWED_46 ,
										MUX_7_1_IN_6 => UNWINDOWED_46 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_23
									);
MUX_REORD_UNIT_24 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_24 ,
										MUX_7_1_IN_1 => UNWINDOWED_24 ,
										MUX_7_1_IN_2 => UNWINDOWED_24 ,
										MUX_7_1_IN_3 => UNWINDOWED_17 ,
										MUX_7_1_IN_4 => UNWINDOWED_17 ,
										MUX_7_1_IN_5 => UNWINDOWED_48 ,
										MUX_7_1_IN_6 => UNWINDOWED_48 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_24
									);
MUX_REORD_UNIT_25 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_25 ,
										MUX_7_1_IN_1 => UNWINDOWED_26 ,
										MUX_7_1_IN_2 => UNWINDOWED_26 ,
										MUX_7_1_IN_3 => UNWINDOWED_19 ,
										MUX_7_1_IN_4 => UNWINDOWED_19 ,
										MUX_7_1_IN_5 => UNWINDOWED_50 ,
										MUX_7_1_IN_6 => UNWINDOWED_50 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_25
									);
MUX_REORD_UNIT_26 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_26 ,
										MUX_7_1_IN_1 => UNWINDOWED_25 ,
										MUX_7_1_IN_2 => UNWINDOWED_28 ,
										MUX_7_1_IN_3 => UNWINDOWED_21 ,
										MUX_7_1_IN_4 => UNWINDOWED_21 ,
										MUX_7_1_IN_5 => UNWINDOWED_52 ,
										MUX_7_1_IN_6 => UNWINDOWED_52 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_26
									);
MUX_REORD_UNIT_27 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_27 ,
										MUX_7_1_IN_1 => UNWINDOWED_27 ,
										MUX_7_1_IN_2 => UNWINDOWED_30 ,
										MUX_7_1_IN_3 => UNWINDOWED_23 ,
										MUX_7_1_IN_4 => UNWINDOWED_23 ,
										MUX_7_1_IN_5 => UNWINDOWED_54 ,
										MUX_7_1_IN_6 => UNWINDOWED_54 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_27
									);
MUX_REORD_UNIT_28 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_28 ,
										MUX_7_1_IN_1 => UNWINDOWED_28 ,
										MUX_7_1_IN_2 => UNWINDOWED_25 ,
										MUX_7_1_IN_3 => UNWINDOWED_25 ,
										MUX_7_1_IN_4 => UNWINDOWED_25 ,
										MUX_7_1_IN_5 => UNWINDOWED_56 ,
										MUX_7_1_IN_6 => UNWINDOWED_56 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_28
									);
MUX_REORD_UNIT_29 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_29 ,
										MUX_7_1_IN_1 => UNWINDOWED_30 ,
										MUX_7_1_IN_2 => UNWINDOWED_27 ,
										MUX_7_1_IN_3 => UNWINDOWED_27 ,
										MUX_7_1_IN_4 => UNWINDOWED_27 ,
										MUX_7_1_IN_5 => UNWINDOWED_58 ,
										MUX_7_1_IN_6 => UNWINDOWED_58 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_29
									);
MUX_REORD_UNIT_30 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_30 ,
										MUX_7_1_IN_1 => UNWINDOWED_29 ,
										MUX_7_1_IN_2 => UNWINDOWED_29 ,
										MUX_7_1_IN_3 => UNWINDOWED_29 ,
										MUX_7_1_IN_4 => UNWINDOWED_29 ,
										MUX_7_1_IN_5 => UNWINDOWED_60 ,
										MUX_7_1_IN_6 => UNWINDOWED_60 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_30
									);
MUX_REORD_UNIT_31 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_31 ,
										MUX_7_1_IN_1 => UNWINDOWED_31 ,
										MUX_7_1_IN_2 => UNWINDOWED_31 ,
										MUX_7_1_IN_3 => UNWINDOWED_31 ,
										MUX_7_1_IN_4 => UNWINDOWED_31 ,
										MUX_7_1_IN_5 => UNWINDOWED_62 ,
										MUX_7_1_IN_6 => UNWINDOWED_62 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_31
									);
MUX_REORD_UNIT_32 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_32 ,
										MUX_7_1_IN_1 => UNWINDOWED_32 ,
										MUX_7_1_IN_2 => UNWINDOWED_32 ,
										MUX_7_1_IN_3 => UNWINDOWED_32 ,
										MUX_7_1_IN_4 => UNWINDOWED_32 ,
										MUX_7_1_IN_5 => UNWINDOWED_1 ,
										MUX_7_1_IN_6 => UNWINDOWED_64 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_32
									);
MUX_REORD_UNIT_33 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_33 ,
										MUX_7_1_IN_1 => UNWINDOWED_34 ,
										MUX_7_1_IN_2 => UNWINDOWED_34 ,
										MUX_7_1_IN_3 => UNWINDOWED_34 ,
										MUX_7_1_IN_4 => UNWINDOWED_34 ,
										MUX_7_1_IN_5 => UNWINDOWED_3 ,
										MUX_7_1_IN_6 => UNWINDOWED_66 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_33
									);
MUX_REORD_UNIT_34 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_34 ,
										MUX_7_1_IN_1 => UNWINDOWED_33 ,
										MUX_7_1_IN_2 => UNWINDOWED_36 ,
										MUX_7_1_IN_3 => UNWINDOWED_36 ,
										MUX_7_1_IN_4 => UNWINDOWED_36 ,
										MUX_7_1_IN_5 => UNWINDOWED_5 ,
										MUX_7_1_IN_6 => UNWINDOWED_68 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_34
									);
MUX_REORD_UNIT_35 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_35 ,
										MUX_7_1_IN_1 => UNWINDOWED_35 ,
										MUX_7_1_IN_2 => UNWINDOWED_38 ,
										MUX_7_1_IN_3 => UNWINDOWED_38 ,
										MUX_7_1_IN_4 => UNWINDOWED_38 ,
										MUX_7_1_IN_5 => UNWINDOWED_7 ,
										MUX_7_1_IN_6 => UNWINDOWED_70 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_35
									);
MUX_REORD_UNIT_36 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_36 ,
										MUX_7_1_IN_1 => UNWINDOWED_36 ,
										MUX_7_1_IN_2 => UNWINDOWED_33 ,
										MUX_7_1_IN_3 => UNWINDOWED_40 ,
										MUX_7_1_IN_4 => UNWINDOWED_40 ,
										MUX_7_1_IN_5 => UNWINDOWED_9 ,
										MUX_7_1_IN_6 => UNWINDOWED_72 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_36
									);
MUX_REORD_UNIT_37 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_37 ,
										MUX_7_1_IN_1 => UNWINDOWED_38 ,
										MUX_7_1_IN_2 => UNWINDOWED_35 ,
										MUX_7_1_IN_3 => UNWINDOWED_42 ,
										MUX_7_1_IN_4 => UNWINDOWED_42 ,
										MUX_7_1_IN_5 => UNWINDOWED_11 ,
										MUX_7_1_IN_6 => UNWINDOWED_74 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_37
									);
MUX_REORD_UNIT_38 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_38 ,
										MUX_7_1_IN_1 => UNWINDOWED_37 ,
										MUX_7_1_IN_2 => UNWINDOWED_37 ,
										MUX_7_1_IN_3 => UNWINDOWED_44 ,
										MUX_7_1_IN_4 => UNWINDOWED_44 ,
										MUX_7_1_IN_5 => UNWINDOWED_13 ,
										MUX_7_1_IN_6 => UNWINDOWED_76 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_38
									);
MUX_REORD_UNIT_39 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_39 ,
										MUX_7_1_IN_1 => UNWINDOWED_39 ,
										MUX_7_1_IN_2 => UNWINDOWED_39 ,
										MUX_7_1_IN_3 => UNWINDOWED_46 ,
										MUX_7_1_IN_4 => UNWINDOWED_46 ,
										MUX_7_1_IN_5 => UNWINDOWED_15 ,
										MUX_7_1_IN_6 => UNWINDOWED_78 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_39
									);
MUX_REORD_UNIT_40 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_40 ,
										MUX_7_1_IN_1 => UNWINDOWED_40 ,
										MUX_7_1_IN_2 => UNWINDOWED_40 ,
										MUX_7_1_IN_3 => UNWINDOWED_33 ,
										MUX_7_1_IN_4 => UNWINDOWED_48 ,
										MUX_7_1_IN_5 => UNWINDOWED_17 ,
										MUX_7_1_IN_6 => UNWINDOWED_80 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_40
									);
MUX_REORD_UNIT_41 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_41 ,
										MUX_7_1_IN_1 => UNWINDOWED_42 ,
										MUX_7_1_IN_2 => UNWINDOWED_42 ,
										MUX_7_1_IN_3 => UNWINDOWED_35 ,
										MUX_7_1_IN_4 => UNWINDOWED_50 ,
										MUX_7_1_IN_5 => UNWINDOWED_19 ,
										MUX_7_1_IN_6 => UNWINDOWED_82 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_41
									);
MUX_REORD_UNIT_42 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_42 ,
										MUX_7_1_IN_1 => UNWINDOWED_41 ,
										MUX_7_1_IN_2 => UNWINDOWED_44 ,
										MUX_7_1_IN_3 => UNWINDOWED_37 ,
										MUX_7_1_IN_4 => UNWINDOWED_52 ,
										MUX_7_1_IN_5 => UNWINDOWED_21 ,
										MUX_7_1_IN_6 => UNWINDOWED_84 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_42
									);
MUX_REORD_UNIT_43 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_43 ,
										MUX_7_1_IN_1 => UNWINDOWED_43 ,
										MUX_7_1_IN_2 => UNWINDOWED_46 ,
										MUX_7_1_IN_3 => UNWINDOWED_39 ,
										MUX_7_1_IN_4 => UNWINDOWED_54 ,
										MUX_7_1_IN_5 => UNWINDOWED_23 ,
										MUX_7_1_IN_6 => UNWINDOWED_86 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_43
									);
MUX_REORD_UNIT_44 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_44 ,
										MUX_7_1_IN_1 => UNWINDOWED_44 ,
										MUX_7_1_IN_2 => UNWINDOWED_41 ,
										MUX_7_1_IN_3 => UNWINDOWED_41 ,
										MUX_7_1_IN_4 => UNWINDOWED_56 ,
										MUX_7_1_IN_5 => UNWINDOWED_25 ,
										MUX_7_1_IN_6 => UNWINDOWED_88 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_44
									);
MUX_REORD_UNIT_45 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_45 ,
										MUX_7_1_IN_1 => UNWINDOWED_46 ,
										MUX_7_1_IN_2 => UNWINDOWED_43 ,
										MUX_7_1_IN_3 => UNWINDOWED_43 ,
										MUX_7_1_IN_4 => UNWINDOWED_58 ,
										MUX_7_1_IN_5 => UNWINDOWED_27 ,
										MUX_7_1_IN_6 => UNWINDOWED_90 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_45
									);
MUX_REORD_UNIT_46 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_46 ,
										MUX_7_1_IN_1 => UNWINDOWED_45 ,
										MUX_7_1_IN_2 => UNWINDOWED_45 ,
										MUX_7_1_IN_3 => UNWINDOWED_45 ,
										MUX_7_1_IN_4 => UNWINDOWED_60 ,
										MUX_7_1_IN_5 => UNWINDOWED_29 ,
										MUX_7_1_IN_6 => UNWINDOWED_92 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_46
									);
MUX_REORD_UNIT_47 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_47 ,
										MUX_7_1_IN_1 => UNWINDOWED_47 ,
										MUX_7_1_IN_2 => UNWINDOWED_47 ,
										MUX_7_1_IN_3 => UNWINDOWED_47 ,
										MUX_7_1_IN_4 => UNWINDOWED_62 ,
										MUX_7_1_IN_5 => UNWINDOWED_31 ,
										MUX_7_1_IN_6 => UNWINDOWED_94 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_47
									);
MUX_REORD_UNIT_48 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_48 ,
										MUX_7_1_IN_1 => UNWINDOWED_48 ,
										MUX_7_1_IN_2 => UNWINDOWED_48 ,
										MUX_7_1_IN_3 => UNWINDOWED_48 ,
										MUX_7_1_IN_4 => UNWINDOWED_33 ,
										MUX_7_1_IN_5 => UNWINDOWED_33 ,
										MUX_7_1_IN_6 => UNWINDOWED_96 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_48
									);
MUX_REORD_UNIT_49 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_49 ,
										MUX_7_1_IN_1 => UNWINDOWED_50 ,
										MUX_7_1_IN_2 => UNWINDOWED_50 ,
										MUX_7_1_IN_3 => UNWINDOWED_50 ,
										MUX_7_1_IN_4 => UNWINDOWED_35 ,
										MUX_7_1_IN_5 => UNWINDOWED_35 ,
										MUX_7_1_IN_6 => UNWINDOWED_98 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_49
									);
MUX_REORD_UNIT_50 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_50 ,
										MUX_7_1_IN_1 => UNWINDOWED_49 ,
										MUX_7_1_IN_2 => UNWINDOWED_52 ,
										MUX_7_1_IN_3 => UNWINDOWED_52 ,
										MUX_7_1_IN_4 => UNWINDOWED_37 ,
										MUX_7_1_IN_5 => UNWINDOWED_37 ,
										MUX_7_1_IN_6 => UNWINDOWED_100 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_50
									);
MUX_REORD_UNIT_51 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_51 ,
										MUX_7_1_IN_1 => UNWINDOWED_51 ,
										MUX_7_1_IN_2 => UNWINDOWED_54 ,
										MUX_7_1_IN_3 => UNWINDOWED_54 ,
										MUX_7_1_IN_4 => UNWINDOWED_39 ,
										MUX_7_1_IN_5 => UNWINDOWED_39 ,
										MUX_7_1_IN_6 => UNWINDOWED_102 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_51
									);
MUX_REORD_UNIT_52 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_52 ,
										MUX_7_1_IN_1 => UNWINDOWED_52 ,
										MUX_7_1_IN_2 => UNWINDOWED_49 ,
										MUX_7_1_IN_3 => UNWINDOWED_56 ,
										MUX_7_1_IN_4 => UNWINDOWED_41 ,
										MUX_7_1_IN_5 => UNWINDOWED_41 ,
										MUX_7_1_IN_6 => UNWINDOWED_104 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_52
									);
MUX_REORD_UNIT_53 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_53 ,
										MUX_7_1_IN_1 => UNWINDOWED_54 ,
										MUX_7_1_IN_2 => UNWINDOWED_51 ,
										MUX_7_1_IN_3 => UNWINDOWED_58 ,
										MUX_7_1_IN_4 => UNWINDOWED_43 ,
										MUX_7_1_IN_5 => UNWINDOWED_43 ,
										MUX_7_1_IN_6 => UNWINDOWED_106 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_53
									);
MUX_REORD_UNIT_54 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_54 ,
										MUX_7_1_IN_1 => UNWINDOWED_53 ,
										MUX_7_1_IN_2 => UNWINDOWED_53 ,
										MUX_7_1_IN_3 => UNWINDOWED_60 ,
										MUX_7_1_IN_4 => UNWINDOWED_45 ,
										MUX_7_1_IN_5 => UNWINDOWED_45 ,
										MUX_7_1_IN_6 => UNWINDOWED_108 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_54
									);
MUX_REORD_UNIT_55 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_55 ,
										MUX_7_1_IN_1 => UNWINDOWED_55 ,
										MUX_7_1_IN_2 => UNWINDOWED_55 ,
										MUX_7_1_IN_3 => UNWINDOWED_62 ,
										MUX_7_1_IN_4 => UNWINDOWED_47 ,
										MUX_7_1_IN_5 => UNWINDOWED_47 ,
										MUX_7_1_IN_6 => UNWINDOWED_110 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_55
									);
MUX_REORD_UNIT_56 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_56 ,
										MUX_7_1_IN_1 => UNWINDOWED_56 ,
										MUX_7_1_IN_2 => UNWINDOWED_56 ,
										MUX_7_1_IN_3 => UNWINDOWED_49 ,
										MUX_7_1_IN_4 => UNWINDOWED_49 ,
										MUX_7_1_IN_5 => UNWINDOWED_49 ,
										MUX_7_1_IN_6 => UNWINDOWED_112 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_56
									);
MUX_REORD_UNIT_57 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_57 ,
										MUX_7_1_IN_1 => UNWINDOWED_58 ,
										MUX_7_1_IN_2 => UNWINDOWED_58 ,
										MUX_7_1_IN_3 => UNWINDOWED_51 ,
										MUX_7_1_IN_4 => UNWINDOWED_51 ,
										MUX_7_1_IN_5 => UNWINDOWED_51 ,
										MUX_7_1_IN_6 => UNWINDOWED_114 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_57
									);
MUX_REORD_UNIT_58 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_58 ,
										MUX_7_1_IN_1 => UNWINDOWED_57 ,
										MUX_7_1_IN_2 => UNWINDOWED_60 ,
										MUX_7_1_IN_3 => UNWINDOWED_53 ,
										MUX_7_1_IN_4 => UNWINDOWED_53 ,
										MUX_7_1_IN_5 => UNWINDOWED_53 ,
										MUX_7_1_IN_6 => UNWINDOWED_116 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_58
									);
MUX_REORD_UNIT_59 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_59 ,
										MUX_7_1_IN_1 => UNWINDOWED_59 ,
										MUX_7_1_IN_2 => UNWINDOWED_62 ,
										MUX_7_1_IN_3 => UNWINDOWED_55 ,
										MUX_7_1_IN_4 => UNWINDOWED_55 ,
										MUX_7_1_IN_5 => UNWINDOWED_55 ,
										MUX_7_1_IN_6 => UNWINDOWED_118 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_59
									);
MUX_REORD_UNIT_60 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_60 ,
										MUX_7_1_IN_1 => UNWINDOWED_60 ,
										MUX_7_1_IN_2 => UNWINDOWED_57 ,
										MUX_7_1_IN_3 => UNWINDOWED_57 ,
										MUX_7_1_IN_4 => UNWINDOWED_57 ,
										MUX_7_1_IN_5 => UNWINDOWED_57 ,
										MUX_7_1_IN_6 => UNWINDOWED_120 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_60
									);
MUX_REORD_UNIT_61 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_61 ,
										MUX_7_1_IN_1 => UNWINDOWED_62 ,
										MUX_7_1_IN_2 => UNWINDOWED_59 ,
										MUX_7_1_IN_3 => UNWINDOWED_59 ,
										MUX_7_1_IN_4 => UNWINDOWED_59 ,
										MUX_7_1_IN_5 => UNWINDOWED_59 ,
										MUX_7_1_IN_6 => UNWINDOWED_122 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_61
									);
MUX_REORD_UNIT_62 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_62 ,
										MUX_7_1_IN_1 => UNWINDOWED_61 ,
										MUX_7_1_IN_2 => UNWINDOWED_61 ,
										MUX_7_1_IN_3 => UNWINDOWED_61 ,
										MUX_7_1_IN_4 => UNWINDOWED_61 ,
										MUX_7_1_IN_5 => UNWINDOWED_61 ,
										MUX_7_1_IN_6 => UNWINDOWED_124 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_62
									);
MUX_REORD_UNIT_63 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_63 ,
										MUX_7_1_IN_1 => UNWINDOWED_63 ,
										MUX_7_1_IN_2 => UNWINDOWED_63 ,
										MUX_7_1_IN_3 => UNWINDOWED_63 ,
										MUX_7_1_IN_4 => UNWINDOWED_63 ,
										MUX_7_1_IN_5 => UNWINDOWED_63 ,
										MUX_7_1_IN_6 => UNWINDOWED_126 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_63
									);
MUX_REORD_UNIT_64 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_64 ,
										MUX_7_1_IN_1 => UNWINDOWED_64 ,
										MUX_7_1_IN_2 => UNWINDOWED_64 ,
										MUX_7_1_IN_3 => UNWINDOWED_64 ,
										MUX_7_1_IN_4 => UNWINDOWED_64 ,
										MUX_7_1_IN_5 => UNWINDOWED_64 ,
										MUX_7_1_IN_6 => UNWINDOWED_1 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_64
									);
MUX_REORD_UNIT_65 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_65 ,
										MUX_7_1_IN_1 => UNWINDOWED_66 ,
										MUX_7_1_IN_2 => UNWINDOWED_66 ,
										MUX_7_1_IN_3 => UNWINDOWED_66 ,
										MUX_7_1_IN_4 => UNWINDOWED_66 ,
										MUX_7_1_IN_5 => UNWINDOWED_66 ,
										MUX_7_1_IN_6 => UNWINDOWED_3 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_65
									);
MUX_REORD_UNIT_66 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_66 ,
										MUX_7_1_IN_1 => UNWINDOWED_65 ,
										MUX_7_1_IN_2 => UNWINDOWED_68 ,
										MUX_7_1_IN_3 => UNWINDOWED_68 ,
										MUX_7_1_IN_4 => UNWINDOWED_68 ,
										MUX_7_1_IN_5 => UNWINDOWED_68 ,
										MUX_7_1_IN_6 => UNWINDOWED_5 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_66
									);
MUX_REORD_UNIT_67 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_67 ,
										MUX_7_1_IN_1 => UNWINDOWED_67 ,
										MUX_7_1_IN_2 => UNWINDOWED_70 ,
										MUX_7_1_IN_3 => UNWINDOWED_70 ,
										MUX_7_1_IN_4 => UNWINDOWED_70 ,
										MUX_7_1_IN_5 => UNWINDOWED_70 ,
										MUX_7_1_IN_6 => UNWINDOWED_7 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_67
									);
MUX_REORD_UNIT_68 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_68 ,
										MUX_7_1_IN_1 => UNWINDOWED_68 ,
										MUX_7_1_IN_2 => UNWINDOWED_65 ,
										MUX_7_1_IN_3 => UNWINDOWED_72 ,
										MUX_7_1_IN_4 => UNWINDOWED_72 ,
										MUX_7_1_IN_5 => UNWINDOWED_72 ,
										MUX_7_1_IN_6 => UNWINDOWED_9 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_68
									);
MUX_REORD_UNIT_69 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_69 ,
										MUX_7_1_IN_1 => UNWINDOWED_70 ,
										MUX_7_1_IN_2 => UNWINDOWED_67 ,
										MUX_7_1_IN_3 => UNWINDOWED_74 ,
										MUX_7_1_IN_4 => UNWINDOWED_74 ,
										MUX_7_1_IN_5 => UNWINDOWED_74 ,
										MUX_7_1_IN_6 => UNWINDOWED_11 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_69
									);
MUX_REORD_UNIT_70 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_70 ,
										MUX_7_1_IN_1 => UNWINDOWED_69 ,
										MUX_7_1_IN_2 => UNWINDOWED_69 ,
										MUX_7_1_IN_3 => UNWINDOWED_76 ,
										MUX_7_1_IN_4 => UNWINDOWED_76 ,
										MUX_7_1_IN_5 => UNWINDOWED_76 ,
										MUX_7_1_IN_6 => UNWINDOWED_13 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_70
									);
MUX_REORD_UNIT_71 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_71 ,
										MUX_7_1_IN_1 => UNWINDOWED_71 ,
										MUX_7_1_IN_2 => UNWINDOWED_71 ,
										MUX_7_1_IN_3 => UNWINDOWED_78 ,
										MUX_7_1_IN_4 => UNWINDOWED_78 ,
										MUX_7_1_IN_5 => UNWINDOWED_78 ,
										MUX_7_1_IN_6 => UNWINDOWED_15 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_71
									);
MUX_REORD_UNIT_72 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_72 ,
										MUX_7_1_IN_1 => UNWINDOWED_72 ,
										MUX_7_1_IN_2 => UNWINDOWED_72 ,
										MUX_7_1_IN_3 => UNWINDOWED_65 ,
										MUX_7_1_IN_4 => UNWINDOWED_80 ,
										MUX_7_1_IN_5 => UNWINDOWED_80 ,
										MUX_7_1_IN_6 => UNWINDOWED_17 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_72
									);
MUX_REORD_UNIT_73 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_73 ,
										MUX_7_1_IN_1 => UNWINDOWED_74 ,
										MUX_7_1_IN_2 => UNWINDOWED_74 ,
										MUX_7_1_IN_3 => UNWINDOWED_67 ,
										MUX_7_1_IN_4 => UNWINDOWED_82 ,
										MUX_7_1_IN_5 => UNWINDOWED_82 ,
										MUX_7_1_IN_6 => UNWINDOWED_19 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_73
									);
MUX_REORD_UNIT_74 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_74 ,
										MUX_7_1_IN_1 => UNWINDOWED_73 ,
										MUX_7_1_IN_2 => UNWINDOWED_76 ,
										MUX_7_1_IN_3 => UNWINDOWED_69 ,
										MUX_7_1_IN_4 => UNWINDOWED_84 ,
										MUX_7_1_IN_5 => UNWINDOWED_84 ,
										MUX_7_1_IN_6 => UNWINDOWED_21 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_74
									);
MUX_REORD_UNIT_75 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_75 ,
										MUX_7_1_IN_1 => UNWINDOWED_75 ,
										MUX_7_1_IN_2 => UNWINDOWED_78 ,
										MUX_7_1_IN_3 => UNWINDOWED_71 ,
										MUX_7_1_IN_4 => UNWINDOWED_86 ,
										MUX_7_1_IN_5 => UNWINDOWED_86 ,
										MUX_7_1_IN_6 => UNWINDOWED_23 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_75
									);
MUX_REORD_UNIT_76 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_76 ,
										MUX_7_1_IN_1 => UNWINDOWED_76 ,
										MUX_7_1_IN_2 => UNWINDOWED_73 ,
										MUX_7_1_IN_3 => UNWINDOWED_73 ,
										MUX_7_1_IN_4 => UNWINDOWED_88 ,
										MUX_7_1_IN_5 => UNWINDOWED_88 ,
										MUX_7_1_IN_6 => UNWINDOWED_25 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_76
									);
MUX_REORD_UNIT_77 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_77 ,
										MUX_7_1_IN_1 => UNWINDOWED_78 ,
										MUX_7_1_IN_2 => UNWINDOWED_75 ,
										MUX_7_1_IN_3 => UNWINDOWED_75 ,
										MUX_7_1_IN_4 => UNWINDOWED_90 ,
										MUX_7_1_IN_5 => UNWINDOWED_90 ,
										MUX_7_1_IN_6 => UNWINDOWED_27 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_77
									);
MUX_REORD_UNIT_78 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_78 ,
										MUX_7_1_IN_1 => UNWINDOWED_77 ,
										MUX_7_1_IN_2 => UNWINDOWED_77 ,
										MUX_7_1_IN_3 => UNWINDOWED_77 ,
										MUX_7_1_IN_4 => UNWINDOWED_92 ,
										MUX_7_1_IN_5 => UNWINDOWED_92 ,
										MUX_7_1_IN_6 => UNWINDOWED_29 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_78
									);
MUX_REORD_UNIT_79 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_79 ,
										MUX_7_1_IN_1 => UNWINDOWED_79 ,
										MUX_7_1_IN_2 => UNWINDOWED_79 ,
										MUX_7_1_IN_3 => UNWINDOWED_79 ,
										MUX_7_1_IN_4 => UNWINDOWED_94 ,
										MUX_7_1_IN_5 => UNWINDOWED_94 ,
										MUX_7_1_IN_6 => UNWINDOWED_31 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_79
									);
MUX_REORD_UNIT_80 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_80 ,
										MUX_7_1_IN_1 => UNWINDOWED_80 ,
										MUX_7_1_IN_2 => UNWINDOWED_80 ,
										MUX_7_1_IN_3 => UNWINDOWED_80 ,
										MUX_7_1_IN_4 => UNWINDOWED_65 ,
										MUX_7_1_IN_5 => UNWINDOWED_96 ,
										MUX_7_1_IN_6 => UNWINDOWED_33 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_80
									);
MUX_REORD_UNIT_81 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_81 ,
										MUX_7_1_IN_1 => UNWINDOWED_82 ,
										MUX_7_1_IN_2 => UNWINDOWED_82 ,
										MUX_7_1_IN_3 => UNWINDOWED_82 ,
										MUX_7_1_IN_4 => UNWINDOWED_67 ,
										MUX_7_1_IN_5 => UNWINDOWED_98 ,
										MUX_7_1_IN_6 => UNWINDOWED_35 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_81
									);
MUX_REORD_UNIT_82 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_82 ,
										MUX_7_1_IN_1 => UNWINDOWED_81 ,
										MUX_7_1_IN_2 => UNWINDOWED_84 ,
										MUX_7_1_IN_3 => UNWINDOWED_84 ,
										MUX_7_1_IN_4 => UNWINDOWED_69 ,
										MUX_7_1_IN_5 => UNWINDOWED_100 ,
										MUX_7_1_IN_6 => UNWINDOWED_37 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_82
									);
MUX_REORD_UNIT_83 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_83 ,
										MUX_7_1_IN_1 => UNWINDOWED_83 ,
										MUX_7_1_IN_2 => UNWINDOWED_86 ,
										MUX_7_1_IN_3 => UNWINDOWED_86 ,
										MUX_7_1_IN_4 => UNWINDOWED_71 ,
										MUX_7_1_IN_5 => UNWINDOWED_102 ,
										MUX_7_1_IN_6 => UNWINDOWED_39 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_83
									);
MUX_REORD_UNIT_84 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_84 ,
										MUX_7_1_IN_1 => UNWINDOWED_84 ,
										MUX_7_1_IN_2 => UNWINDOWED_81 ,
										MUX_7_1_IN_3 => UNWINDOWED_88 ,
										MUX_7_1_IN_4 => UNWINDOWED_73 ,
										MUX_7_1_IN_5 => UNWINDOWED_104 ,
										MUX_7_1_IN_6 => UNWINDOWED_41 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_84
									);
MUX_REORD_UNIT_85 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_85 ,
										MUX_7_1_IN_1 => UNWINDOWED_86 ,
										MUX_7_1_IN_2 => UNWINDOWED_83 ,
										MUX_7_1_IN_3 => UNWINDOWED_90 ,
										MUX_7_1_IN_4 => UNWINDOWED_75 ,
										MUX_7_1_IN_5 => UNWINDOWED_106 ,
										MUX_7_1_IN_6 => UNWINDOWED_43 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_85
									);
MUX_REORD_UNIT_86 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_86 ,
										MUX_7_1_IN_1 => UNWINDOWED_85 ,
										MUX_7_1_IN_2 => UNWINDOWED_85 ,
										MUX_7_1_IN_3 => UNWINDOWED_92 ,
										MUX_7_1_IN_4 => UNWINDOWED_77 ,
										MUX_7_1_IN_5 => UNWINDOWED_108 ,
										MUX_7_1_IN_6 => UNWINDOWED_45 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_86
									);
MUX_REORD_UNIT_87 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_87 ,
										MUX_7_1_IN_1 => UNWINDOWED_87 ,
										MUX_7_1_IN_2 => UNWINDOWED_87 ,
										MUX_7_1_IN_3 => UNWINDOWED_94 ,
										MUX_7_1_IN_4 => UNWINDOWED_79 ,
										MUX_7_1_IN_5 => UNWINDOWED_110 ,
										MUX_7_1_IN_6 => UNWINDOWED_47 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_87
									);
MUX_REORD_UNIT_88 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_88 ,
										MUX_7_1_IN_1 => UNWINDOWED_88 ,
										MUX_7_1_IN_2 => UNWINDOWED_88 ,
										MUX_7_1_IN_3 => UNWINDOWED_81 ,
										MUX_7_1_IN_4 => UNWINDOWED_81 ,
										MUX_7_1_IN_5 => UNWINDOWED_112 ,
										MUX_7_1_IN_6 => UNWINDOWED_49 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_88
									);
MUX_REORD_UNIT_89 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_89 ,
										MUX_7_1_IN_1 => UNWINDOWED_90 ,
										MUX_7_1_IN_2 => UNWINDOWED_90 ,
										MUX_7_1_IN_3 => UNWINDOWED_83 ,
										MUX_7_1_IN_4 => UNWINDOWED_83 ,
										MUX_7_1_IN_5 => UNWINDOWED_114 ,
										MUX_7_1_IN_6 => UNWINDOWED_51 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_89
									);
MUX_REORD_UNIT_90 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_90 ,
										MUX_7_1_IN_1 => UNWINDOWED_89 ,
										MUX_7_1_IN_2 => UNWINDOWED_92 ,
										MUX_7_1_IN_3 => UNWINDOWED_85 ,
										MUX_7_1_IN_4 => UNWINDOWED_85 ,
										MUX_7_1_IN_5 => UNWINDOWED_116 ,
										MUX_7_1_IN_6 => UNWINDOWED_53 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_90
									);
MUX_REORD_UNIT_91 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_91 ,
										MUX_7_1_IN_1 => UNWINDOWED_91 ,
										MUX_7_1_IN_2 => UNWINDOWED_94 ,
										MUX_7_1_IN_3 => UNWINDOWED_87 ,
										MUX_7_1_IN_4 => UNWINDOWED_87 ,
										MUX_7_1_IN_5 => UNWINDOWED_118 ,
										MUX_7_1_IN_6 => UNWINDOWED_55 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_91
									);
MUX_REORD_UNIT_92 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_92 ,
										MUX_7_1_IN_1 => UNWINDOWED_92 ,
										MUX_7_1_IN_2 => UNWINDOWED_89 ,
										MUX_7_1_IN_3 => UNWINDOWED_89 ,
										MUX_7_1_IN_4 => UNWINDOWED_89 ,
										MUX_7_1_IN_5 => UNWINDOWED_120 ,
										MUX_7_1_IN_6 => UNWINDOWED_57 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_92
									);
MUX_REORD_UNIT_93 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_93 ,
										MUX_7_1_IN_1 => UNWINDOWED_94 ,
										MUX_7_1_IN_2 => UNWINDOWED_91 ,
										MUX_7_1_IN_3 => UNWINDOWED_91 ,
										MUX_7_1_IN_4 => UNWINDOWED_91 ,
										MUX_7_1_IN_5 => UNWINDOWED_122 ,
										MUX_7_1_IN_6 => UNWINDOWED_59 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_93
									);
MUX_REORD_UNIT_94 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_94 ,
										MUX_7_1_IN_1 => UNWINDOWED_93 ,
										MUX_7_1_IN_2 => UNWINDOWED_93 ,
										MUX_7_1_IN_3 => UNWINDOWED_93 ,
										MUX_7_1_IN_4 => UNWINDOWED_93 ,
										MUX_7_1_IN_5 => UNWINDOWED_124 ,
										MUX_7_1_IN_6 => UNWINDOWED_61 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_94
									);
MUX_REORD_UNIT_95 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_95 ,
										MUX_7_1_IN_1 => UNWINDOWED_95 ,
										MUX_7_1_IN_2 => UNWINDOWED_95 ,
										MUX_7_1_IN_3 => UNWINDOWED_95 ,
										MUX_7_1_IN_4 => UNWINDOWED_95 ,
										MUX_7_1_IN_5 => UNWINDOWED_126 ,
										MUX_7_1_IN_6 => UNWINDOWED_63 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_95
									);
MUX_REORD_UNIT_96 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_96 ,
										MUX_7_1_IN_1 => UNWINDOWED_96 ,
										MUX_7_1_IN_2 => UNWINDOWED_96 ,
										MUX_7_1_IN_3 => UNWINDOWED_96 ,
										MUX_7_1_IN_4 => UNWINDOWED_96 ,
										MUX_7_1_IN_5 => UNWINDOWED_65 ,
										MUX_7_1_IN_6 => UNWINDOWED_65 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_96
									);
MUX_REORD_UNIT_97 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_97 ,
										MUX_7_1_IN_1 => UNWINDOWED_98 ,
										MUX_7_1_IN_2 => UNWINDOWED_98 ,
										MUX_7_1_IN_3 => UNWINDOWED_98 ,
										MUX_7_1_IN_4 => UNWINDOWED_98 ,
										MUX_7_1_IN_5 => UNWINDOWED_67 ,
										MUX_7_1_IN_6 => UNWINDOWED_67 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_97
									);
MUX_REORD_UNIT_98 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_98 ,
										MUX_7_1_IN_1 => UNWINDOWED_97 ,
										MUX_7_1_IN_2 => UNWINDOWED_100 ,
										MUX_7_1_IN_3 => UNWINDOWED_100 ,
										MUX_7_1_IN_4 => UNWINDOWED_100 ,
										MUX_7_1_IN_5 => UNWINDOWED_69 ,
										MUX_7_1_IN_6 => UNWINDOWED_69 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_98
									);
MUX_REORD_UNIT_99 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_99 ,
										MUX_7_1_IN_1 => UNWINDOWED_99 ,
										MUX_7_1_IN_2 => UNWINDOWED_102 ,
										MUX_7_1_IN_3 => UNWINDOWED_102 ,
										MUX_7_1_IN_4 => UNWINDOWED_102 ,
										MUX_7_1_IN_5 => UNWINDOWED_71 ,
										MUX_7_1_IN_6 => UNWINDOWED_71 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_99
									);
MUX_REORD_UNIT_100 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_100 ,
										MUX_7_1_IN_1 => UNWINDOWED_100 ,
										MUX_7_1_IN_2 => UNWINDOWED_97 ,
										MUX_7_1_IN_3 => UNWINDOWED_104 ,
										MUX_7_1_IN_4 => UNWINDOWED_104 ,
										MUX_7_1_IN_5 => UNWINDOWED_73 ,
										MUX_7_1_IN_6 => UNWINDOWED_73 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_100
									);
MUX_REORD_UNIT_101 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_101 ,
										MUX_7_1_IN_1 => UNWINDOWED_102 ,
										MUX_7_1_IN_2 => UNWINDOWED_99 ,
										MUX_7_1_IN_3 => UNWINDOWED_106 ,
										MUX_7_1_IN_4 => UNWINDOWED_106 ,
										MUX_7_1_IN_5 => UNWINDOWED_75 ,
										MUX_7_1_IN_6 => UNWINDOWED_75 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_101
									);
MUX_REORD_UNIT_102 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_102 ,
										MUX_7_1_IN_1 => UNWINDOWED_101 ,
										MUX_7_1_IN_2 => UNWINDOWED_101 ,
										MUX_7_1_IN_3 => UNWINDOWED_108 ,
										MUX_7_1_IN_4 => UNWINDOWED_108 ,
										MUX_7_1_IN_5 => UNWINDOWED_77 ,
										MUX_7_1_IN_6 => UNWINDOWED_77 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_102
									);
MUX_REORD_UNIT_103 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_103 ,
										MUX_7_1_IN_1 => UNWINDOWED_103 ,
										MUX_7_1_IN_2 => UNWINDOWED_103 ,
										MUX_7_1_IN_3 => UNWINDOWED_110 ,
										MUX_7_1_IN_4 => UNWINDOWED_110 ,
										MUX_7_1_IN_5 => UNWINDOWED_79 ,
										MUX_7_1_IN_6 => UNWINDOWED_79 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_103
									);
MUX_REORD_UNIT_104 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_104 ,
										MUX_7_1_IN_1 => UNWINDOWED_104 ,
										MUX_7_1_IN_2 => UNWINDOWED_104 ,
										MUX_7_1_IN_3 => UNWINDOWED_97 ,
										MUX_7_1_IN_4 => UNWINDOWED_112 ,
										MUX_7_1_IN_5 => UNWINDOWED_81 ,
										MUX_7_1_IN_6 => UNWINDOWED_81 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_104
									);
MUX_REORD_UNIT_105 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_105 ,
										MUX_7_1_IN_1 => UNWINDOWED_106 ,
										MUX_7_1_IN_2 => UNWINDOWED_106 ,
										MUX_7_1_IN_3 => UNWINDOWED_99 ,
										MUX_7_1_IN_4 => UNWINDOWED_114 ,
										MUX_7_1_IN_5 => UNWINDOWED_83 ,
										MUX_7_1_IN_6 => UNWINDOWED_83 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_105
									);
MUX_REORD_UNIT_106 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_106 ,
										MUX_7_1_IN_1 => UNWINDOWED_105 ,
										MUX_7_1_IN_2 => UNWINDOWED_108 ,
										MUX_7_1_IN_3 => UNWINDOWED_101 ,
										MUX_7_1_IN_4 => UNWINDOWED_116 ,
										MUX_7_1_IN_5 => UNWINDOWED_85 ,
										MUX_7_1_IN_6 => UNWINDOWED_85 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_106
									);
MUX_REORD_UNIT_107 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_107 ,
										MUX_7_1_IN_1 => UNWINDOWED_107 ,
										MUX_7_1_IN_2 => UNWINDOWED_110 ,
										MUX_7_1_IN_3 => UNWINDOWED_103 ,
										MUX_7_1_IN_4 => UNWINDOWED_118 ,
										MUX_7_1_IN_5 => UNWINDOWED_87 ,
										MUX_7_1_IN_6 => UNWINDOWED_87 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_107
									);
MUX_REORD_UNIT_108 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_108 ,
										MUX_7_1_IN_1 => UNWINDOWED_108 ,
										MUX_7_1_IN_2 => UNWINDOWED_105 ,
										MUX_7_1_IN_3 => UNWINDOWED_105 ,
										MUX_7_1_IN_4 => UNWINDOWED_120 ,
										MUX_7_1_IN_5 => UNWINDOWED_89 ,
										MUX_7_1_IN_6 => UNWINDOWED_89 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_108
									);
MUX_REORD_UNIT_109 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_109 ,
										MUX_7_1_IN_1 => UNWINDOWED_110 ,
										MUX_7_1_IN_2 => UNWINDOWED_107 ,
										MUX_7_1_IN_3 => UNWINDOWED_107 ,
										MUX_7_1_IN_4 => UNWINDOWED_122 ,
										MUX_7_1_IN_5 => UNWINDOWED_91 ,
										MUX_7_1_IN_6 => UNWINDOWED_91 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_109
									);
MUX_REORD_UNIT_110 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_110 ,
										MUX_7_1_IN_1 => UNWINDOWED_109 ,
										MUX_7_1_IN_2 => UNWINDOWED_109 ,
										MUX_7_1_IN_3 => UNWINDOWED_109 ,
										MUX_7_1_IN_4 => UNWINDOWED_124 ,
										MUX_7_1_IN_5 => UNWINDOWED_93 ,
										MUX_7_1_IN_6 => UNWINDOWED_93 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_110
									);
MUX_REORD_UNIT_111 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_111 ,
										MUX_7_1_IN_1 => UNWINDOWED_111 ,
										MUX_7_1_IN_2 => UNWINDOWED_111 ,
										MUX_7_1_IN_3 => UNWINDOWED_111 ,
										MUX_7_1_IN_4 => UNWINDOWED_126 ,
										MUX_7_1_IN_5 => UNWINDOWED_95 ,
										MUX_7_1_IN_6 => UNWINDOWED_95 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_111
									);
MUX_REORD_UNIT_112 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_112 ,
										MUX_7_1_IN_1 => UNWINDOWED_112 ,
										MUX_7_1_IN_2 => UNWINDOWED_112 ,
										MUX_7_1_IN_3 => UNWINDOWED_112 ,
										MUX_7_1_IN_4 => UNWINDOWED_97 ,
										MUX_7_1_IN_5 => UNWINDOWED_97 ,
										MUX_7_1_IN_6 => UNWINDOWED_97 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_112
									);
MUX_REORD_UNIT_113 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_113 ,
										MUX_7_1_IN_1 => UNWINDOWED_114 ,
										MUX_7_1_IN_2 => UNWINDOWED_114 ,
										MUX_7_1_IN_3 => UNWINDOWED_114 ,
										MUX_7_1_IN_4 => UNWINDOWED_99 ,
										MUX_7_1_IN_5 => UNWINDOWED_99 ,
										MUX_7_1_IN_6 => UNWINDOWED_99 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_113
									);
MUX_REORD_UNIT_114 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_114 ,
										MUX_7_1_IN_1 => UNWINDOWED_113 ,
										MUX_7_1_IN_2 => UNWINDOWED_116 ,
										MUX_7_1_IN_3 => UNWINDOWED_116 ,
										MUX_7_1_IN_4 => UNWINDOWED_101 ,
										MUX_7_1_IN_5 => UNWINDOWED_101 ,
										MUX_7_1_IN_6 => UNWINDOWED_101 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_114
									);
MUX_REORD_UNIT_115 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_115 ,
										MUX_7_1_IN_1 => UNWINDOWED_115 ,
										MUX_7_1_IN_2 => UNWINDOWED_118 ,
										MUX_7_1_IN_3 => UNWINDOWED_118 ,
										MUX_7_1_IN_4 => UNWINDOWED_103 ,
										MUX_7_1_IN_5 => UNWINDOWED_103 ,
										MUX_7_1_IN_6 => UNWINDOWED_103 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_115
									);
MUX_REORD_UNIT_116 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_116 ,
										MUX_7_1_IN_1 => UNWINDOWED_116 ,
										MUX_7_1_IN_2 => UNWINDOWED_113 ,
										MUX_7_1_IN_3 => UNWINDOWED_120 ,
										MUX_7_1_IN_4 => UNWINDOWED_105 ,
										MUX_7_1_IN_5 => UNWINDOWED_105 ,
										MUX_7_1_IN_6 => UNWINDOWED_105 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_116
									);
MUX_REORD_UNIT_117 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_117 ,
										MUX_7_1_IN_1 => UNWINDOWED_118 ,
										MUX_7_1_IN_2 => UNWINDOWED_115 ,
										MUX_7_1_IN_3 => UNWINDOWED_122 ,
										MUX_7_1_IN_4 => UNWINDOWED_107 ,
										MUX_7_1_IN_5 => UNWINDOWED_107 ,
										MUX_7_1_IN_6 => UNWINDOWED_107 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_117
									);
MUX_REORD_UNIT_118 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_118 ,
										MUX_7_1_IN_1 => UNWINDOWED_117 ,
										MUX_7_1_IN_2 => UNWINDOWED_117 ,
										MUX_7_1_IN_3 => UNWINDOWED_124 ,
										MUX_7_1_IN_4 => UNWINDOWED_109 ,
										MUX_7_1_IN_5 => UNWINDOWED_109 ,
										MUX_7_1_IN_6 => UNWINDOWED_109 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_118
									);
MUX_REORD_UNIT_119 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_119 ,
										MUX_7_1_IN_1 => UNWINDOWED_119 ,
										MUX_7_1_IN_2 => UNWINDOWED_119 ,
										MUX_7_1_IN_3 => UNWINDOWED_126 ,
										MUX_7_1_IN_4 => UNWINDOWED_111 ,
										MUX_7_1_IN_5 => UNWINDOWED_111 ,
										MUX_7_1_IN_6 => UNWINDOWED_111 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_119
									);
MUX_REORD_UNIT_120 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_120 ,
										MUX_7_1_IN_1 => UNWINDOWED_120 ,
										MUX_7_1_IN_2 => UNWINDOWED_120 ,
										MUX_7_1_IN_3 => UNWINDOWED_113 ,
										MUX_7_1_IN_4 => UNWINDOWED_113 ,
										MUX_7_1_IN_5 => UNWINDOWED_113 ,
										MUX_7_1_IN_6 => UNWINDOWED_113 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_120
									);
MUX_REORD_UNIT_121 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_121 ,
										MUX_7_1_IN_1 => UNWINDOWED_122 ,
										MUX_7_1_IN_2 => UNWINDOWED_122 ,
										MUX_7_1_IN_3 => UNWINDOWED_115 ,
										MUX_7_1_IN_4 => UNWINDOWED_115 ,
										MUX_7_1_IN_5 => UNWINDOWED_115 ,
										MUX_7_1_IN_6 => UNWINDOWED_115 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_121
									);
MUX_REORD_UNIT_122 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_122 ,
										MUX_7_1_IN_1 => UNWINDOWED_121 ,
										MUX_7_1_IN_2 => UNWINDOWED_124 ,
										MUX_7_1_IN_3 => UNWINDOWED_117 ,
										MUX_7_1_IN_4 => UNWINDOWED_117 ,
										MUX_7_1_IN_5 => UNWINDOWED_117 ,
										MUX_7_1_IN_6 => UNWINDOWED_117 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_122
									);
MUX_REORD_UNIT_123 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_123 ,
										MUX_7_1_IN_1 => UNWINDOWED_123 ,
										MUX_7_1_IN_2 => UNWINDOWED_126 ,
										MUX_7_1_IN_3 => UNWINDOWED_119 ,
										MUX_7_1_IN_4 => UNWINDOWED_119 ,
										MUX_7_1_IN_5 => UNWINDOWED_119 ,
										MUX_7_1_IN_6 => UNWINDOWED_119 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_123
									);
MUX_REORD_UNIT_124 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_124 ,
										MUX_7_1_IN_1 => UNWINDOWED_124 ,
										MUX_7_1_IN_2 => UNWINDOWED_121 ,
										MUX_7_1_IN_3 => UNWINDOWED_121 ,
										MUX_7_1_IN_4 => UNWINDOWED_121 ,
										MUX_7_1_IN_5 => UNWINDOWED_121 ,
										MUX_7_1_IN_6 => UNWINDOWED_121 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_124
									);
MUX_REORD_UNIT_125 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_125 ,
										MUX_7_1_IN_1 => UNWINDOWED_126 ,
										MUX_7_1_IN_2 => UNWINDOWED_123 ,
										MUX_7_1_IN_3 => UNWINDOWED_123 ,
										MUX_7_1_IN_4 => UNWINDOWED_123 ,
										MUX_7_1_IN_5 => UNWINDOWED_123 ,
										MUX_7_1_IN_6 => UNWINDOWED_123 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_125
									);
MUX_REORD_UNIT_126 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_126 ,
										MUX_7_1_IN_1 => UNWINDOWED_125 ,
										MUX_7_1_IN_2 => UNWINDOWED_125 ,
										MUX_7_1_IN_3 => UNWINDOWED_125 ,
										MUX_7_1_IN_4 => UNWINDOWED_125 ,
										MUX_7_1_IN_5 => UNWINDOWED_125 ,
										MUX_7_1_IN_6 => UNWINDOWED_125 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_126
									);
MUX_REORD_UNIT_127 : multiplexer_7_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_7_1_IN_0 => UNWINDOWED_127 ,
										MUX_7_1_IN_1 => UNWINDOWED_127 ,
										MUX_7_1_IN_2 => UNWINDOWED_127 ,
										MUX_7_1_IN_3 => UNWINDOWED_127 ,
										MUX_7_1_IN_4 => UNWINDOWED_127 ,
										MUX_7_1_IN_5 => UNWINDOWED_127 ,
										MUX_7_1_IN_6 => UNWINDOWED_127 ,
				                    			MUX_7_1_IN_SEL => QEP_N_7_W_5_S_0_IN_QTGT ,
										MUX_7_1_OUT_RES => TO_STATE_REG_127
									);

MUX_OUTPUT_SELECTION : multiplexer_128_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_128_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_128_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_128_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_128_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_128_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_128_1_IN_5 => FROM_STATE_REG_5 ,
										MUX_128_1_IN_6 => FROM_STATE_REG_6 ,
										MUX_128_1_IN_7 => FROM_STATE_REG_7 ,
										MUX_128_1_IN_8 => FROM_STATE_REG_8 ,
										MUX_128_1_IN_9 => FROM_STATE_REG_9 ,
										MUX_128_1_IN_10 => FROM_STATE_REG_10 ,
										MUX_128_1_IN_11 => FROM_STATE_REG_11 ,
										MUX_128_1_IN_12 => FROM_STATE_REG_12 ,
										MUX_128_1_IN_13 => FROM_STATE_REG_13 ,
										MUX_128_1_IN_14 => FROM_STATE_REG_14 ,
										MUX_128_1_IN_15 => FROM_STATE_REG_15 ,
										MUX_128_1_IN_16 => FROM_STATE_REG_16 ,
										MUX_128_1_IN_17 => FROM_STATE_REG_17 ,
										MUX_128_1_IN_18 => FROM_STATE_REG_18 ,
										MUX_128_1_IN_19 => FROM_STATE_REG_19 ,
										MUX_128_1_IN_20 => FROM_STATE_REG_20 ,
										MUX_128_1_IN_21 => FROM_STATE_REG_21 ,
										MUX_128_1_IN_22 => FROM_STATE_REG_22 ,
										MUX_128_1_IN_23 => FROM_STATE_REG_23 ,
										MUX_128_1_IN_24 => FROM_STATE_REG_24 ,
										MUX_128_1_IN_25 => FROM_STATE_REG_25 ,
										MUX_128_1_IN_26 => FROM_STATE_REG_26 ,
										MUX_128_1_IN_27 => FROM_STATE_REG_27 ,
										MUX_128_1_IN_28 => FROM_STATE_REG_28 ,
										MUX_128_1_IN_29 => FROM_STATE_REG_29 ,
										MUX_128_1_IN_30 => FROM_STATE_REG_30 ,
										MUX_128_1_IN_31 => FROM_STATE_REG_31 ,
										MUX_128_1_IN_32 => FROM_STATE_REG_32 ,
										MUX_128_1_IN_33 => FROM_STATE_REG_33 ,
										MUX_128_1_IN_34 => FROM_STATE_REG_34 ,
										MUX_128_1_IN_35 => FROM_STATE_REG_35 ,
										MUX_128_1_IN_36 => FROM_STATE_REG_36 ,
										MUX_128_1_IN_37 => FROM_STATE_REG_37 ,
										MUX_128_1_IN_38 => FROM_STATE_REG_38 ,
										MUX_128_1_IN_39 => FROM_STATE_REG_39 ,
										MUX_128_1_IN_40 => FROM_STATE_REG_40 ,
										MUX_128_1_IN_41 => FROM_STATE_REG_41 ,
										MUX_128_1_IN_42 => FROM_STATE_REG_42 ,
										MUX_128_1_IN_43 => FROM_STATE_REG_43 ,
										MUX_128_1_IN_44 => FROM_STATE_REG_44 ,
										MUX_128_1_IN_45 => FROM_STATE_REG_45 ,
										MUX_128_1_IN_46 => FROM_STATE_REG_46 ,
										MUX_128_1_IN_47 => FROM_STATE_REG_47 ,
										MUX_128_1_IN_48 => FROM_STATE_REG_48 ,
										MUX_128_1_IN_49 => FROM_STATE_REG_49 ,
										MUX_128_1_IN_50 => FROM_STATE_REG_50 ,
										MUX_128_1_IN_51 => FROM_STATE_REG_51 ,
										MUX_128_1_IN_52 => FROM_STATE_REG_52 ,
										MUX_128_1_IN_53 => FROM_STATE_REG_53 ,
										MUX_128_1_IN_54 => FROM_STATE_REG_54 ,
										MUX_128_1_IN_55 => FROM_STATE_REG_55 ,
										MUX_128_1_IN_56 => FROM_STATE_REG_56 ,
										MUX_128_1_IN_57 => FROM_STATE_REG_57 ,
										MUX_128_1_IN_58 => FROM_STATE_REG_58 ,
										MUX_128_1_IN_59 => FROM_STATE_REG_59 ,
										MUX_128_1_IN_60 => FROM_STATE_REG_60 ,
										MUX_128_1_IN_61 => FROM_STATE_REG_61 ,
										MUX_128_1_IN_62 => FROM_STATE_REG_62 ,
										MUX_128_1_IN_63 => FROM_STATE_REG_63 ,
										MUX_128_1_IN_64 => FROM_STATE_REG_64 ,
										MUX_128_1_IN_65 => FROM_STATE_REG_65 ,
										MUX_128_1_IN_66 => FROM_STATE_REG_66 ,
										MUX_128_1_IN_67 => FROM_STATE_REG_67 ,
										MUX_128_1_IN_68 => FROM_STATE_REG_68 ,
										MUX_128_1_IN_69 => FROM_STATE_REG_69 ,
										MUX_128_1_IN_70 => FROM_STATE_REG_70 ,
										MUX_128_1_IN_71 => FROM_STATE_REG_71 ,
										MUX_128_1_IN_72 => FROM_STATE_REG_72 ,
										MUX_128_1_IN_73 => FROM_STATE_REG_73 ,
										MUX_128_1_IN_74 => FROM_STATE_REG_74 ,
										MUX_128_1_IN_75 => FROM_STATE_REG_75 ,
										MUX_128_1_IN_76 => FROM_STATE_REG_76 ,
										MUX_128_1_IN_77 => FROM_STATE_REG_77 ,
										MUX_128_1_IN_78 => FROM_STATE_REG_78 ,
										MUX_128_1_IN_79 => FROM_STATE_REG_79 ,
										MUX_128_1_IN_80 => FROM_STATE_REG_80 ,
										MUX_128_1_IN_81 => FROM_STATE_REG_81 ,
										MUX_128_1_IN_82 => FROM_STATE_REG_82 ,
										MUX_128_1_IN_83 => FROM_STATE_REG_83 ,
										MUX_128_1_IN_84 => FROM_STATE_REG_84 ,
										MUX_128_1_IN_85 => FROM_STATE_REG_85 ,
										MUX_128_1_IN_86 => FROM_STATE_REG_86 ,
										MUX_128_1_IN_87 => FROM_STATE_REG_87 ,
										MUX_128_1_IN_88 => FROM_STATE_REG_88 ,
										MUX_128_1_IN_89 => FROM_STATE_REG_89 ,
										MUX_128_1_IN_90 => FROM_STATE_REG_90 ,
										MUX_128_1_IN_91 => FROM_STATE_REG_91 ,
										MUX_128_1_IN_92 => FROM_STATE_REG_92 ,
										MUX_128_1_IN_93 => FROM_STATE_REG_93 ,
										MUX_128_1_IN_94 => FROM_STATE_REG_94 ,
										MUX_128_1_IN_95 => FROM_STATE_REG_95 ,
										MUX_128_1_IN_96 => FROM_STATE_REG_96 ,
										MUX_128_1_IN_97 => FROM_STATE_REG_97 ,
										MUX_128_1_IN_98 => FROM_STATE_REG_98 ,
										MUX_128_1_IN_99 => FROM_STATE_REG_99 ,
										MUX_128_1_IN_100 => FROM_STATE_REG_100 ,
										MUX_128_1_IN_101 => FROM_STATE_REG_101 ,
										MUX_128_1_IN_102 => FROM_STATE_REG_102 ,
										MUX_128_1_IN_103 => FROM_STATE_REG_103 ,
										MUX_128_1_IN_104 => FROM_STATE_REG_104 ,
										MUX_128_1_IN_105 => FROM_STATE_REG_105 ,
										MUX_128_1_IN_106 => FROM_STATE_REG_106 ,
										MUX_128_1_IN_107 => FROM_STATE_REG_107 ,
										MUX_128_1_IN_108 => FROM_STATE_REG_108 ,
										MUX_128_1_IN_109 => FROM_STATE_REG_109 ,
										MUX_128_1_IN_110 => FROM_STATE_REG_110 ,
										MUX_128_1_IN_111 => FROM_STATE_REG_111 ,
										MUX_128_1_IN_112 => FROM_STATE_REG_112 ,
										MUX_128_1_IN_113 => FROM_STATE_REG_113 ,
										MUX_128_1_IN_114 => FROM_STATE_REG_114 ,
										MUX_128_1_IN_115 => FROM_STATE_REG_115 ,
										MUX_128_1_IN_116 => FROM_STATE_REG_116 ,
										MUX_128_1_IN_117 => FROM_STATE_REG_117 ,
										MUX_128_1_IN_118 => FROM_STATE_REG_118 ,
										MUX_128_1_IN_119 => FROM_STATE_REG_119 ,
										MUX_128_1_IN_120 => FROM_STATE_REG_120 ,
										MUX_128_1_IN_121 => FROM_STATE_REG_121 ,
										MUX_128_1_IN_122 => FROM_STATE_REG_122 ,
										MUX_128_1_IN_123 => FROM_STATE_REG_123 ,
										MUX_128_1_IN_124 => FROM_STATE_REG_124 ,
										MUX_128_1_IN_125 => FROM_STATE_REG_125 ,
										MUX_128_1_IN_126 => FROM_STATE_REG_126 ,
										MUX_128_1_IN_127 => FROM_STATE_REG_127 ,
				                    			MUX_128_1_IN_SEL => QEP_N_7_W_5_S_0_IN_OUT_STATE_SEL ,
										MUX_128_1_OUT_RES => SELECTED_OUTPUT
									);
MUX_REAL_IMAG_SELECTION : multiplexer_2_1 GENERIC MAP (K => K)
									PORT MAP (
										MUX_2_1_IN_0 => SELECTED_OUTPUT((2*K-1) DOWNTO K),
										MUX_2_1_IN_1 => SELECTED_OUTPUT((K-1) DOWNTO 0),
				                    			MUX_2_1_IN_SEL => QEP_N_7_W_5_S_0_IN_REAL_IMAG_SEL ,
										MUX_2_1_OUT_RES => QEP_N_7_W_5_S_0_OUT_DATA
									);

END generated;