LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY rot_rom IS 	
	PORT(
		ROT_ROM_IN_ADD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		ROT_ROM_OUT : OUT STD_LOGIC_VECTOR (41 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF rot_rom IS

BEGIN

--Output signal follows the pattern
-- |DONE|NEXT_ADD|CTRL_INST|
-- |  1 |  5     |   36    |
--CTRL_INST is divided as follows
-- |PIPE|LD|OBI|OBR|OAI|OAR|S1A|S1B|S2A|S2B|M12A|M1B|M2B|SUB|SAVED|
-- | 3  |3 | 3 | 2 | 2 | 2 | 3 | 2 | 2 | 2 |  1 | 3 | 3 | 2 |  3  |

-- 					   DONE  NEXT_ADD    PIPE    LD      OBI    OBR    OAI    OAR     S1A    S1B    S2A    S2B   M12A    M1B     M2B   SUB     SAVED
-- 						1	     5         3      3       3       2      2      2      3      2 	 2      2     1       3       3     2        3  
	ROT_ROM_OUT <= 
						'0' & "00100" & "001" & "000" & "000" & "00" & "00" & "00" & "000" & "00" & "00" & "00" & '0' & "000" & "011" & "00" & "000"	
						 WHEN ROT_ROM_IN_ADD = "00000" ELSE		--RX_I
						
						'0' & "00101" & "001" & "000" & "000" & "00" & "00" & "00" & "000" & "00" & "00" & "00" & '0' & "000" & "010" & "00" & "000"	
						 WHEN ROT_ROM_IN_ADD = "00001" ELSE		--RY_I
						
						'0' & "00110" & "001" & "000" & "000" & "00" & "00" & "00" & "000" & "00" & "00" & "00" & '0' & "000" & "001" & "00" & "000"	
						 WHEN ROT_ROM_IN_ADD = "00010" ELSE		--RZ_I
						
						'0' & "00111" & "001" & "000" & "000" & "00" & "00" & "00" & "000" & "00" & "00" & "00" & '0' & "010" & "011" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "00011" ELSE		--U1_I
						
						'0' & "01000" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "00100" ELSE		--RX_II
						
						'0' & "01001" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "00101" ELSE		--RY_II
						
						'0' & "01010" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "00110" ELSE		--RZ_II
						
						'0' & "01011" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "00111" ELSE		--U1_II
						
						'0' & "01100" & "001" & "001" & "000" & "00" & "00" & "10" & "011" & "10" & "00" & "00" & '0' & "001" & "010" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "01000" ELSE		--RX_III
						
						'0' & "01101" & "001" & "001" & "000" & "00" & "00" & "10" & "011" & "10" & "00" & "00" & '0' & "001" & "011" & "01" & "000"
						 WHEN ROT_ROM_IN_ADD = "01001" ELSE		--RY_III
												
						'0' & "01110" & "001" & "001" & "000" & "00" & "00" & "10" & "011" & "10" & "00" & "00" & '0' & "001" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "01010" ELSE		--RZ_III
												
						'0' & "01111" & "001" & "100" & "000" & "10" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "011" & "010" & "01" & "000"
						 WHEN ROT_ROM_IN_ADD = "01011" ELSE		--U1_III
												
						'0' & "10000" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "01100" ELSE		--RX_IV
						
						'0' & "10001" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "01101" ELSE		--RY_IV
						
						'0' & "10010" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "01110" ELSE		--RZ_IV
						
						'0' & "10011" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "01111" ELSE		--U1_IV
						
						'0' & "10100" & "001" & "010" & "000" & "00" & "10" & "00" & "011" & "10" & "00" & "00" & '0' & "010" & "001" & "01" & "000"	
						 WHEN ROT_ROM_IN_ADD = "10000" ELSE		--RX_V
						
						'0' & "11001" & "001" & "010" & "000" & "00" & "10" & "00" & "011" & "10" & "00" & "00" & '0' & "010" & "000" & "01" & "000"	
						 WHEN ROT_ROM_IN_ADD = "10001" ELSE		--RY_V
						
						'0' & "11010" & "001" & "010" & "000" & "00" & "10" & "00" & "011" & "10" & "00" & "00" & '0' & "010" & "011" & "01" & "000"	
						 WHEN ROT_ROM_IN_ADD = "10010" ELSE		--RZ_V
						
						'1' & "00000" & "000" & "000" & "010" & "00" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "000" & "000" & "00" & "100"
						 WHEN ROT_ROM_IN_ADD = "10011" ELSE		--U1_V
						
						'0' & "10101" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "10100" ELSE		--RX_VI
						
						'0' & "10110" & "001" & "100" & "000" & "10" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "011" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "10101" ELSE		--RX_VII
						
						'0' & "10111" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "10110" ELSE		--RX_VIII
						
						'1' & "00000" & "000" & "000" & "010" & "00" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "000" & "000" & "01" & "111"
						 WHEN ROT_ROM_IN_ADD = "10111" ELSE		--RX_IX
						
						'1' & "00000" & "000" & "000" & "010" & "00" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "000" & "000" & "00" & "111"
						 WHEN ROT_ROM_IN_ADD = "11000" ELSE		--RZ_IX
						
						'0' & "11011" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "11001" ELSE		--RY_VI
												
						'0' & "11100" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "11010" ELSE		--RZ_VI
												
						'0' & "11101" & "001" & "100" & "000" & "10" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "011" & "001" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "11011" ELSE		--RY_VII
												
						'0' & "11110" & "001" & "100" & "000" & "10" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "011" & "010" & "01" & "000"
						 WHEN ROT_ROM_IN_ADD = "11100" ELSE		--RZ_VII
						
						'0' & "11111" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "11101" ELSE		--RY_VIII
						
						'0' & "11000" & "100" & "000" & "000" & "00" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN ROT_ROM_IN_ADD = "11110" ELSE		--RZ_VIII
						
						'1' & "00000" & "000" & "000" & "010" & "00" & "00" & "00" & "011" & "10" & "00" & "00" & '0' & "000" & "000" & "00" & "111"
						 WHEN ROT_ROM_IN_ADD = "11111" ELSE		--RY_IX
						
						
						(OTHERS => '0');

END behavioral;