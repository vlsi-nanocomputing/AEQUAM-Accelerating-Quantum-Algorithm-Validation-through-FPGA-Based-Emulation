library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_1024_1 IS 
	GENERIC (K : INTEGER := 40);
	PORT (
		MUX_1024_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_32 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_33 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_34 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_35 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_36 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_37 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_38 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_39 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_40 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_41 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_42 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_43 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_44 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_45 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_46 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_47 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_48 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_49 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_50 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_51 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_52 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_53 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_54 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_55 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_56 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_57 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_58 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_59 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_60 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_61 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_62 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_63 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_64 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_65 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_66 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_67 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_68 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_69 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_70 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_71 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_72 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_73 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_74 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_75 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_76 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_77 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_78 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_79 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_80 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_81 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_82 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_83 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_84 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_85 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_86 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_87 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_88 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_89 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_90 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_91 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_92 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_93 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_94 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_95 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_96 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_97 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_98 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_99 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_100 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_101 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_102 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_103 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_104 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_105 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_106 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_107 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_108 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_109 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_110 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_111 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_112 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_113 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_114 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_115 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_116 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_117 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_118 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_119 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_120 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_121 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_122 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_123 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_124 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_125 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_126 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_127 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_128 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_129 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_130 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_131 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_132 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_133 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_134 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_135 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_136 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_137 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_138 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_139 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_140 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_141 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_142 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_143 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_144 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_145 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_146 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_147 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_148 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_149 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_150 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_151 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_152 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_153 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_154 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_155 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_156 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_157 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_158 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_159 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_160 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_161 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_162 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_163 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_164 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_165 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_166 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_167 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_168 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_169 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_170 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_171 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_172 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_173 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_174 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_175 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_176 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_177 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_178 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_179 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_180 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_181 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_182 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_183 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_184 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_185 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_186 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_187 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_188 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_189 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_190 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_191 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_192 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_193 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_194 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_195 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_196 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_197 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_198 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_199 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_200 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_201 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_202 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_203 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_204 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_205 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_206 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_207 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_208 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_209 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_210 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_211 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_212 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_213 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_214 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_215 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_216 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_217 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_218 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_219 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_220 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_221 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_222 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_223 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_224 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_225 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_226 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_227 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_228 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_229 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_230 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_231 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_232 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_233 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_234 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_235 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_236 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_237 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_238 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_239 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_240 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_241 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_242 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_243 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_244 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_245 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_246 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_247 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_248 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_249 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_250 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_251 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_252 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_253 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_254 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_255 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_256 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_257 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_258 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_259 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_260 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_261 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_262 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_263 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_264 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_265 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_266 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_267 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_268 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_269 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_270 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_271 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_272 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_273 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_274 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_275 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_276 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_277 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_278 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_279 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_280 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_281 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_282 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_283 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_284 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_285 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_286 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_287 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_288 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_289 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_290 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_291 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_292 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_293 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_294 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_295 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_296 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_297 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_298 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_299 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_300 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_301 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_302 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_303 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_304 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_305 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_306 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_307 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_308 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_309 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_310 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_311 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_312 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_313 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_314 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_315 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_316 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_317 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_318 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_319 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_320 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_321 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_322 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_323 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_324 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_325 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_326 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_327 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_328 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_329 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_330 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_331 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_332 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_333 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_334 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_335 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_336 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_337 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_338 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_339 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_340 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_341 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_342 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_343 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_344 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_345 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_346 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_347 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_348 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_349 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_350 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_351 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_352 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_353 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_354 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_355 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_356 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_357 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_358 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_359 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_360 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_361 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_362 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_363 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_364 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_365 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_366 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_367 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_368 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_369 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_370 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_371 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_372 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_373 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_374 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_375 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_376 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_377 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_378 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_379 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_380 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_381 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_382 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_383 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_384 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_385 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_386 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_387 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_388 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_389 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_390 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_391 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_392 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_393 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_394 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_395 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_396 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_397 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_398 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_399 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_400 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_401 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_402 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_403 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_404 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_405 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_406 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_407 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_408 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_409 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_410 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_411 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_412 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_413 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_414 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_415 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_416 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_417 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_418 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_419 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_420 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_421 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_422 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_423 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_424 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_425 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_426 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_427 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_428 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_429 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_430 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_431 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_432 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_433 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_434 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_435 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_436 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_437 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_438 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_439 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_440 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_441 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_442 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_443 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_444 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_445 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_446 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_447 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_448 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_449 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_450 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_451 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_452 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_453 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_454 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_455 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_456 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_457 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_458 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_459 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_460 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_461 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_462 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_463 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_464 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_465 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_466 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_467 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_468 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_469 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_470 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_471 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_472 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_473 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_474 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_475 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_476 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_477 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_478 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_479 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_480 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_481 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_482 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_483 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_484 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_485 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_486 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_487 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_488 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_489 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_490 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_491 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_492 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_493 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_494 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_495 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_496 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_497 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_498 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_499 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_500 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_501 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_502 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_503 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_504 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_505 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_506 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_507 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_508 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_509 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_510 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_511 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_512 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_513 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_514 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_515 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_516 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_517 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_518 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_519 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_520 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_521 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_522 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_523 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_524 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_525 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_526 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_527 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_528 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_529 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_530 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_531 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_532 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_533 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_534 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_535 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_536 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_537 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_538 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_539 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_540 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_541 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_542 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_543 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_544 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_545 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_546 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_547 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_548 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_549 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_550 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_551 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_552 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_553 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_554 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_555 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_556 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_557 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_558 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_559 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_560 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_561 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_562 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_563 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_564 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_565 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_566 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_567 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_568 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_569 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_570 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_571 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_572 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_573 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_574 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_575 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_576 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_577 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_578 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_579 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_580 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_581 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_582 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_583 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_584 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_585 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_586 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_587 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_588 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_589 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_590 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_591 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_592 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_593 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_594 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_595 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_596 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_597 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_598 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_599 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_600 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_601 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_602 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_603 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_604 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_605 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_606 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_607 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_608 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_609 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_610 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_611 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_612 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_613 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_614 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_615 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_616 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_617 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_618 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_619 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_620 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_621 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_622 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_623 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_624 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_625 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_626 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_627 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_628 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_629 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_630 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_631 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_632 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_633 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_634 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_635 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_636 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_637 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_638 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_639 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_640 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_641 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_642 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_643 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_644 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_645 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_646 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_647 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_648 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_649 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_650 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_651 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_652 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_653 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_654 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_655 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_656 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_657 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_658 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_659 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_660 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_661 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_662 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_663 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_664 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_665 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_666 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_667 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_668 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_669 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_670 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_671 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_672 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_673 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_674 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_675 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_676 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_677 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_678 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_679 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_680 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_681 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_682 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_683 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_684 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_685 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_686 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_687 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_688 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_689 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_690 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_691 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_692 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_693 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_694 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_695 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_696 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_697 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_698 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_699 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_700 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_701 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_702 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_703 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_704 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_705 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_706 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_707 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_708 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_709 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_710 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_711 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_712 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_713 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_714 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_715 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_716 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_717 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_718 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_719 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_720 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_721 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_722 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_723 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_724 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_725 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_726 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_727 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_728 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_729 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_730 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_731 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_732 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_733 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_734 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_735 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_736 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_737 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_738 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_739 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_740 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_741 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_742 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_743 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_744 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_745 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_746 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_747 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_748 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_749 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_750 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_751 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_752 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_753 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_754 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_755 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_756 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_757 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_758 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_759 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_760 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_761 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_762 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_763 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_764 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_765 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_766 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_767 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_768 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_769 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_770 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_771 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_772 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_773 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_774 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_775 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_776 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_777 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_778 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_779 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_780 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_781 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_782 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_783 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_784 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_785 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_786 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_787 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_788 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_789 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_790 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_791 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_792 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_793 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_794 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_795 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_796 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_797 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_798 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_799 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_800 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_801 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_802 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_803 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_804 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_805 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_806 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_807 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_808 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_809 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_810 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_811 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_812 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_813 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_814 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_815 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_816 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_817 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_818 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_819 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_820 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_821 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_822 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_823 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_824 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_825 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_826 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_827 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_828 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_829 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_830 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_831 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_832 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_833 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_834 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_835 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_836 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_837 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_838 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_839 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_840 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_841 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_842 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_843 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_844 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_845 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_846 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_847 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_848 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_849 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_850 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_851 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_852 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_853 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_854 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_855 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_856 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_857 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_858 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_859 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_860 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_861 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_862 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_863 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_864 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_865 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_866 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_867 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_868 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_869 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_870 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_871 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_872 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_873 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_874 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_875 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_876 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_877 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_878 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_879 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_880 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_881 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_882 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_883 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_884 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_885 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_886 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_887 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_888 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_889 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_890 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_891 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_892 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_893 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_894 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_895 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_896 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_897 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_898 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_899 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_900 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_901 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_902 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_903 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_904 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_905 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_906 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_907 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_908 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_909 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_910 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_911 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_912 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_913 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_914 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_915 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_916 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_917 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_918 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_919 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_920 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_921 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_922 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_923 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_924 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_925 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_926 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_927 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_928 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_929 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_930 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_931 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_932 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_933 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_934 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_935 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_936 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_937 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_938 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_939 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_940 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_941 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_942 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_943 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_944 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_945 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_946 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_947 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_948 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_949 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_950 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_951 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_952 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_953 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_954 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_955 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_956 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_957 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_958 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_959 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_960 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_961 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_962 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_963 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_964 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_965 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_966 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_967 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_968 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_969 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_970 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_971 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_972 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_973 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_974 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_975 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_976 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_977 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_978 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_979 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_980 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_981 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_982 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_983 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_984 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_985 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_986 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_987 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_988 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_989 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_990 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_991 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_992 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_993 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_994 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_995 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_996 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_997 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_998 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_999 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1000 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1001 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1002 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1003 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1004 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1005 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1006 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1007 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1008 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1009 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1010 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1011 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1012 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1013 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1014 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1015 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1016 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1017 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1018 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1019 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1020 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1021 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1022 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_1023 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1024_1_IN_SEL : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		MUX_1024_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_1024_1 IS

BEGIN

	MUX_1024_1_OUT_RES <= 
				MUX_1024_1_IN_0 WHEN MUX_1024_1_IN_SEL = "0000000000" ELSE
				MUX_1024_1_IN_1 WHEN MUX_1024_1_IN_SEL = "0000000001" ELSE
				MUX_1024_1_IN_2 WHEN MUX_1024_1_IN_SEL = "0000000010" ELSE
				MUX_1024_1_IN_3 WHEN MUX_1024_1_IN_SEL = "0000000011" ELSE
				MUX_1024_1_IN_4 WHEN MUX_1024_1_IN_SEL = "0000000100" ELSE
				MUX_1024_1_IN_5 WHEN MUX_1024_1_IN_SEL = "0000000101" ELSE
				MUX_1024_1_IN_6 WHEN MUX_1024_1_IN_SEL = "0000000110" ELSE
				MUX_1024_1_IN_7 WHEN MUX_1024_1_IN_SEL = "0000000111" ELSE
				MUX_1024_1_IN_8 WHEN MUX_1024_1_IN_SEL = "0000001000" ELSE
				MUX_1024_1_IN_9 WHEN MUX_1024_1_IN_SEL = "0000001001" ELSE
				MUX_1024_1_IN_10 WHEN MUX_1024_1_IN_SEL = "0000001010" ELSE
				MUX_1024_1_IN_11 WHEN MUX_1024_1_IN_SEL = "0000001011" ELSE
				MUX_1024_1_IN_12 WHEN MUX_1024_1_IN_SEL = "0000001100" ELSE
				MUX_1024_1_IN_13 WHEN MUX_1024_1_IN_SEL = "0000001101" ELSE
				MUX_1024_1_IN_14 WHEN MUX_1024_1_IN_SEL = "0000001110" ELSE
				MUX_1024_1_IN_15 WHEN MUX_1024_1_IN_SEL = "0000001111" ELSE
				MUX_1024_1_IN_16 WHEN MUX_1024_1_IN_SEL = "0000010000" ELSE
				MUX_1024_1_IN_17 WHEN MUX_1024_1_IN_SEL = "0000010001" ELSE
				MUX_1024_1_IN_18 WHEN MUX_1024_1_IN_SEL = "0000010010" ELSE
				MUX_1024_1_IN_19 WHEN MUX_1024_1_IN_SEL = "0000010011" ELSE
				MUX_1024_1_IN_20 WHEN MUX_1024_1_IN_SEL = "0000010100" ELSE
				MUX_1024_1_IN_21 WHEN MUX_1024_1_IN_SEL = "0000010101" ELSE
				MUX_1024_1_IN_22 WHEN MUX_1024_1_IN_SEL = "0000010110" ELSE
				MUX_1024_1_IN_23 WHEN MUX_1024_1_IN_SEL = "0000010111" ELSE
				MUX_1024_1_IN_24 WHEN MUX_1024_1_IN_SEL = "0000011000" ELSE
				MUX_1024_1_IN_25 WHEN MUX_1024_1_IN_SEL = "0000011001" ELSE
				MUX_1024_1_IN_26 WHEN MUX_1024_1_IN_SEL = "0000011010" ELSE
				MUX_1024_1_IN_27 WHEN MUX_1024_1_IN_SEL = "0000011011" ELSE
				MUX_1024_1_IN_28 WHEN MUX_1024_1_IN_SEL = "0000011100" ELSE
				MUX_1024_1_IN_29 WHEN MUX_1024_1_IN_SEL = "0000011101" ELSE
				MUX_1024_1_IN_30 WHEN MUX_1024_1_IN_SEL = "0000011110" ELSE
				MUX_1024_1_IN_31 WHEN MUX_1024_1_IN_SEL = "0000011111" ELSE
				MUX_1024_1_IN_32 WHEN MUX_1024_1_IN_SEL = "0000100000" ELSE
				MUX_1024_1_IN_33 WHEN MUX_1024_1_IN_SEL = "0000100001" ELSE
				MUX_1024_1_IN_34 WHEN MUX_1024_1_IN_SEL = "0000100010" ELSE
				MUX_1024_1_IN_35 WHEN MUX_1024_1_IN_SEL = "0000100011" ELSE
				MUX_1024_1_IN_36 WHEN MUX_1024_1_IN_SEL = "0000100100" ELSE
				MUX_1024_1_IN_37 WHEN MUX_1024_1_IN_SEL = "0000100101" ELSE
				MUX_1024_1_IN_38 WHEN MUX_1024_1_IN_SEL = "0000100110" ELSE
				MUX_1024_1_IN_39 WHEN MUX_1024_1_IN_SEL = "0000100111" ELSE
				MUX_1024_1_IN_40 WHEN MUX_1024_1_IN_SEL = "0000101000" ELSE
				MUX_1024_1_IN_41 WHEN MUX_1024_1_IN_SEL = "0000101001" ELSE
				MUX_1024_1_IN_42 WHEN MUX_1024_1_IN_SEL = "0000101010" ELSE
				MUX_1024_1_IN_43 WHEN MUX_1024_1_IN_SEL = "0000101011" ELSE
				MUX_1024_1_IN_44 WHEN MUX_1024_1_IN_SEL = "0000101100" ELSE
				MUX_1024_1_IN_45 WHEN MUX_1024_1_IN_SEL = "0000101101" ELSE
				MUX_1024_1_IN_46 WHEN MUX_1024_1_IN_SEL = "0000101110" ELSE
				MUX_1024_1_IN_47 WHEN MUX_1024_1_IN_SEL = "0000101111" ELSE
				MUX_1024_1_IN_48 WHEN MUX_1024_1_IN_SEL = "0000110000" ELSE
				MUX_1024_1_IN_49 WHEN MUX_1024_1_IN_SEL = "0000110001" ELSE
				MUX_1024_1_IN_50 WHEN MUX_1024_1_IN_SEL = "0000110010" ELSE
				MUX_1024_1_IN_51 WHEN MUX_1024_1_IN_SEL = "0000110011" ELSE
				MUX_1024_1_IN_52 WHEN MUX_1024_1_IN_SEL = "0000110100" ELSE
				MUX_1024_1_IN_53 WHEN MUX_1024_1_IN_SEL = "0000110101" ELSE
				MUX_1024_1_IN_54 WHEN MUX_1024_1_IN_SEL = "0000110110" ELSE
				MUX_1024_1_IN_55 WHEN MUX_1024_1_IN_SEL = "0000110111" ELSE
				MUX_1024_1_IN_56 WHEN MUX_1024_1_IN_SEL = "0000111000" ELSE
				MUX_1024_1_IN_57 WHEN MUX_1024_1_IN_SEL = "0000111001" ELSE
				MUX_1024_1_IN_58 WHEN MUX_1024_1_IN_SEL = "0000111010" ELSE
				MUX_1024_1_IN_59 WHEN MUX_1024_1_IN_SEL = "0000111011" ELSE
				MUX_1024_1_IN_60 WHEN MUX_1024_1_IN_SEL = "0000111100" ELSE
				MUX_1024_1_IN_61 WHEN MUX_1024_1_IN_SEL = "0000111101" ELSE
				MUX_1024_1_IN_62 WHEN MUX_1024_1_IN_SEL = "0000111110" ELSE
				MUX_1024_1_IN_63 WHEN MUX_1024_1_IN_SEL = "0000111111" ELSE
				MUX_1024_1_IN_64 WHEN MUX_1024_1_IN_SEL = "0001000000" ELSE
				MUX_1024_1_IN_65 WHEN MUX_1024_1_IN_SEL = "0001000001" ELSE
				MUX_1024_1_IN_66 WHEN MUX_1024_1_IN_SEL = "0001000010" ELSE
				MUX_1024_1_IN_67 WHEN MUX_1024_1_IN_SEL = "0001000011" ELSE
				MUX_1024_1_IN_68 WHEN MUX_1024_1_IN_SEL = "0001000100" ELSE
				MUX_1024_1_IN_69 WHEN MUX_1024_1_IN_SEL = "0001000101" ELSE
				MUX_1024_1_IN_70 WHEN MUX_1024_1_IN_SEL = "0001000110" ELSE
				MUX_1024_1_IN_71 WHEN MUX_1024_1_IN_SEL = "0001000111" ELSE
				MUX_1024_1_IN_72 WHEN MUX_1024_1_IN_SEL = "0001001000" ELSE
				MUX_1024_1_IN_73 WHEN MUX_1024_1_IN_SEL = "0001001001" ELSE
				MUX_1024_1_IN_74 WHEN MUX_1024_1_IN_SEL = "0001001010" ELSE
				MUX_1024_1_IN_75 WHEN MUX_1024_1_IN_SEL = "0001001011" ELSE
				MUX_1024_1_IN_76 WHEN MUX_1024_1_IN_SEL = "0001001100" ELSE
				MUX_1024_1_IN_77 WHEN MUX_1024_1_IN_SEL = "0001001101" ELSE
				MUX_1024_1_IN_78 WHEN MUX_1024_1_IN_SEL = "0001001110" ELSE
				MUX_1024_1_IN_79 WHEN MUX_1024_1_IN_SEL = "0001001111" ELSE
				MUX_1024_1_IN_80 WHEN MUX_1024_1_IN_SEL = "0001010000" ELSE
				MUX_1024_1_IN_81 WHEN MUX_1024_1_IN_SEL = "0001010001" ELSE
				MUX_1024_1_IN_82 WHEN MUX_1024_1_IN_SEL = "0001010010" ELSE
				MUX_1024_1_IN_83 WHEN MUX_1024_1_IN_SEL = "0001010011" ELSE
				MUX_1024_1_IN_84 WHEN MUX_1024_1_IN_SEL = "0001010100" ELSE
				MUX_1024_1_IN_85 WHEN MUX_1024_1_IN_SEL = "0001010101" ELSE
				MUX_1024_1_IN_86 WHEN MUX_1024_1_IN_SEL = "0001010110" ELSE
				MUX_1024_1_IN_87 WHEN MUX_1024_1_IN_SEL = "0001010111" ELSE
				MUX_1024_1_IN_88 WHEN MUX_1024_1_IN_SEL = "0001011000" ELSE
				MUX_1024_1_IN_89 WHEN MUX_1024_1_IN_SEL = "0001011001" ELSE
				MUX_1024_1_IN_90 WHEN MUX_1024_1_IN_SEL = "0001011010" ELSE
				MUX_1024_1_IN_91 WHEN MUX_1024_1_IN_SEL = "0001011011" ELSE
				MUX_1024_1_IN_92 WHEN MUX_1024_1_IN_SEL = "0001011100" ELSE
				MUX_1024_1_IN_93 WHEN MUX_1024_1_IN_SEL = "0001011101" ELSE
				MUX_1024_1_IN_94 WHEN MUX_1024_1_IN_SEL = "0001011110" ELSE
				MUX_1024_1_IN_95 WHEN MUX_1024_1_IN_SEL = "0001011111" ELSE
				MUX_1024_1_IN_96 WHEN MUX_1024_1_IN_SEL = "0001100000" ELSE
				MUX_1024_1_IN_97 WHEN MUX_1024_1_IN_SEL = "0001100001" ELSE
				MUX_1024_1_IN_98 WHEN MUX_1024_1_IN_SEL = "0001100010" ELSE
				MUX_1024_1_IN_99 WHEN MUX_1024_1_IN_SEL = "0001100011" ELSE
				MUX_1024_1_IN_100 WHEN MUX_1024_1_IN_SEL = "0001100100" ELSE
				MUX_1024_1_IN_101 WHEN MUX_1024_1_IN_SEL = "0001100101" ELSE
				MUX_1024_1_IN_102 WHEN MUX_1024_1_IN_SEL = "0001100110" ELSE
				MUX_1024_1_IN_103 WHEN MUX_1024_1_IN_SEL = "0001100111" ELSE
				MUX_1024_1_IN_104 WHEN MUX_1024_1_IN_SEL = "0001101000" ELSE
				MUX_1024_1_IN_105 WHEN MUX_1024_1_IN_SEL = "0001101001" ELSE
				MUX_1024_1_IN_106 WHEN MUX_1024_1_IN_SEL = "0001101010" ELSE
				MUX_1024_1_IN_107 WHEN MUX_1024_1_IN_SEL = "0001101011" ELSE
				MUX_1024_1_IN_108 WHEN MUX_1024_1_IN_SEL = "0001101100" ELSE
				MUX_1024_1_IN_109 WHEN MUX_1024_1_IN_SEL = "0001101101" ELSE
				MUX_1024_1_IN_110 WHEN MUX_1024_1_IN_SEL = "0001101110" ELSE
				MUX_1024_1_IN_111 WHEN MUX_1024_1_IN_SEL = "0001101111" ELSE
				MUX_1024_1_IN_112 WHEN MUX_1024_1_IN_SEL = "0001110000" ELSE
				MUX_1024_1_IN_113 WHEN MUX_1024_1_IN_SEL = "0001110001" ELSE
				MUX_1024_1_IN_114 WHEN MUX_1024_1_IN_SEL = "0001110010" ELSE
				MUX_1024_1_IN_115 WHEN MUX_1024_1_IN_SEL = "0001110011" ELSE
				MUX_1024_1_IN_116 WHEN MUX_1024_1_IN_SEL = "0001110100" ELSE
				MUX_1024_1_IN_117 WHEN MUX_1024_1_IN_SEL = "0001110101" ELSE
				MUX_1024_1_IN_118 WHEN MUX_1024_1_IN_SEL = "0001110110" ELSE
				MUX_1024_1_IN_119 WHEN MUX_1024_1_IN_SEL = "0001110111" ELSE
				MUX_1024_1_IN_120 WHEN MUX_1024_1_IN_SEL = "0001111000" ELSE
				MUX_1024_1_IN_121 WHEN MUX_1024_1_IN_SEL = "0001111001" ELSE
				MUX_1024_1_IN_122 WHEN MUX_1024_1_IN_SEL = "0001111010" ELSE
				MUX_1024_1_IN_123 WHEN MUX_1024_1_IN_SEL = "0001111011" ELSE
				MUX_1024_1_IN_124 WHEN MUX_1024_1_IN_SEL = "0001111100" ELSE
				MUX_1024_1_IN_125 WHEN MUX_1024_1_IN_SEL = "0001111101" ELSE
				MUX_1024_1_IN_126 WHEN MUX_1024_1_IN_SEL = "0001111110" ELSE
				MUX_1024_1_IN_127 WHEN MUX_1024_1_IN_SEL = "0001111111" ELSE
				MUX_1024_1_IN_128 WHEN MUX_1024_1_IN_SEL = "0010000000" ELSE
				MUX_1024_1_IN_129 WHEN MUX_1024_1_IN_SEL = "0010000001" ELSE
				MUX_1024_1_IN_130 WHEN MUX_1024_1_IN_SEL = "0010000010" ELSE
				MUX_1024_1_IN_131 WHEN MUX_1024_1_IN_SEL = "0010000011" ELSE
				MUX_1024_1_IN_132 WHEN MUX_1024_1_IN_SEL = "0010000100" ELSE
				MUX_1024_1_IN_133 WHEN MUX_1024_1_IN_SEL = "0010000101" ELSE
				MUX_1024_1_IN_134 WHEN MUX_1024_1_IN_SEL = "0010000110" ELSE
				MUX_1024_1_IN_135 WHEN MUX_1024_1_IN_SEL = "0010000111" ELSE
				MUX_1024_1_IN_136 WHEN MUX_1024_1_IN_SEL = "0010001000" ELSE
				MUX_1024_1_IN_137 WHEN MUX_1024_1_IN_SEL = "0010001001" ELSE
				MUX_1024_1_IN_138 WHEN MUX_1024_1_IN_SEL = "0010001010" ELSE
				MUX_1024_1_IN_139 WHEN MUX_1024_1_IN_SEL = "0010001011" ELSE
				MUX_1024_1_IN_140 WHEN MUX_1024_1_IN_SEL = "0010001100" ELSE
				MUX_1024_1_IN_141 WHEN MUX_1024_1_IN_SEL = "0010001101" ELSE
				MUX_1024_1_IN_142 WHEN MUX_1024_1_IN_SEL = "0010001110" ELSE
				MUX_1024_1_IN_143 WHEN MUX_1024_1_IN_SEL = "0010001111" ELSE
				MUX_1024_1_IN_144 WHEN MUX_1024_1_IN_SEL = "0010010000" ELSE
				MUX_1024_1_IN_145 WHEN MUX_1024_1_IN_SEL = "0010010001" ELSE
				MUX_1024_1_IN_146 WHEN MUX_1024_1_IN_SEL = "0010010010" ELSE
				MUX_1024_1_IN_147 WHEN MUX_1024_1_IN_SEL = "0010010011" ELSE
				MUX_1024_1_IN_148 WHEN MUX_1024_1_IN_SEL = "0010010100" ELSE
				MUX_1024_1_IN_149 WHEN MUX_1024_1_IN_SEL = "0010010101" ELSE
				MUX_1024_1_IN_150 WHEN MUX_1024_1_IN_SEL = "0010010110" ELSE
				MUX_1024_1_IN_151 WHEN MUX_1024_1_IN_SEL = "0010010111" ELSE
				MUX_1024_1_IN_152 WHEN MUX_1024_1_IN_SEL = "0010011000" ELSE
				MUX_1024_1_IN_153 WHEN MUX_1024_1_IN_SEL = "0010011001" ELSE
				MUX_1024_1_IN_154 WHEN MUX_1024_1_IN_SEL = "0010011010" ELSE
				MUX_1024_1_IN_155 WHEN MUX_1024_1_IN_SEL = "0010011011" ELSE
				MUX_1024_1_IN_156 WHEN MUX_1024_1_IN_SEL = "0010011100" ELSE
				MUX_1024_1_IN_157 WHEN MUX_1024_1_IN_SEL = "0010011101" ELSE
				MUX_1024_1_IN_158 WHEN MUX_1024_1_IN_SEL = "0010011110" ELSE
				MUX_1024_1_IN_159 WHEN MUX_1024_1_IN_SEL = "0010011111" ELSE
				MUX_1024_1_IN_160 WHEN MUX_1024_1_IN_SEL = "0010100000" ELSE
				MUX_1024_1_IN_161 WHEN MUX_1024_1_IN_SEL = "0010100001" ELSE
				MUX_1024_1_IN_162 WHEN MUX_1024_1_IN_SEL = "0010100010" ELSE
				MUX_1024_1_IN_163 WHEN MUX_1024_1_IN_SEL = "0010100011" ELSE
				MUX_1024_1_IN_164 WHEN MUX_1024_1_IN_SEL = "0010100100" ELSE
				MUX_1024_1_IN_165 WHEN MUX_1024_1_IN_SEL = "0010100101" ELSE
				MUX_1024_1_IN_166 WHEN MUX_1024_1_IN_SEL = "0010100110" ELSE
				MUX_1024_1_IN_167 WHEN MUX_1024_1_IN_SEL = "0010100111" ELSE
				MUX_1024_1_IN_168 WHEN MUX_1024_1_IN_SEL = "0010101000" ELSE
				MUX_1024_1_IN_169 WHEN MUX_1024_1_IN_SEL = "0010101001" ELSE
				MUX_1024_1_IN_170 WHEN MUX_1024_1_IN_SEL = "0010101010" ELSE
				MUX_1024_1_IN_171 WHEN MUX_1024_1_IN_SEL = "0010101011" ELSE
				MUX_1024_1_IN_172 WHEN MUX_1024_1_IN_SEL = "0010101100" ELSE
				MUX_1024_1_IN_173 WHEN MUX_1024_1_IN_SEL = "0010101101" ELSE
				MUX_1024_1_IN_174 WHEN MUX_1024_1_IN_SEL = "0010101110" ELSE
				MUX_1024_1_IN_175 WHEN MUX_1024_1_IN_SEL = "0010101111" ELSE
				MUX_1024_1_IN_176 WHEN MUX_1024_1_IN_SEL = "0010110000" ELSE
				MUX_1024_1_IN_177 WHEN MUX_1024_1_IN_SEL = "0010110001" ELSE
				MUX_1024_1_IN_178 WHEN MUX_1024_1_IN_SEL = "0010110010" ELSE
				MUX_1024_1_IN_179 WHEN MUX_1024_1_IN_SEL = "0010110011" ELSE
				MUX_1024_1_IN_180 WHEN MUX_1024_1_IN_SEL = "0010110100" ELSE
				MUX_1024_1_IN_181 WHEN MUX_1024_1_IN_SEL = "0010110101" ELSE
				MUX_1024_1_IN_182 WHEN MUX_1024_1_IN_SEL = "0010110110" ELSE
				MUX_1024_1_IN_183 WHEN MUX_1024_1_IN_SEL = "0010110111" ELSE
				MUX_1024_1_IN_184 WHEN MUX_1024_1_IN_SEL = "0010111000" ELSE
				MUX_1024_1_IN_185 WHEN MUX_1024_1_IN_SEL = "0010111001" ELSE
				MUX_1024_1_IN_186 WHEN MUX_1024_1_IN_SEL = "0010111010" ELSE
				MUX_1024_1_IN_187 WHEN MUX_1024_1_IN_SEL = "0010111011" ELSE
				MUX_1024_1_IN_188 WHEN MUX_1024_1_IN_SEL = "0010111100" ELSE
				MUX_1024_1_IN_189 WHEN MUX_1024_1_IN_SEL = "0010111101" ELSE
				MUX_1024_1_IN_190 WHEN MUX_1024_1_IN_SEL = "0010111110" ELSE
				MUX_1024_1_IN_191 WHEN MUX_1024_1_IN_SEL = "0010111111" ELSE
				MUX_1024_1_IN_192 WHEN MUX_1024_1_IN_SEL = "0011000000" ELSE
				MUX_1024_1_IN_193 WHEN MUX_1024_1_IN_SEL = "0011000001" ELSE
				MUX_1024_1_IN_194 WHEN MUX_1024_1_IN_SEL = "0011000010" ELSE
				MUX_1024_1_IN_195 WHEN MUX_1024_1_IN_SEL = "0011000011" ELSE
				MUX_1024_1_IN_196 WHEN MUX_1024_1_IN_SEL = "0011000100" ELSE
				MUX_1024_1_IN_197 WHEN MUX_1024_1_IN_SEL = "0011000101" ELSE
				MUX_1024_1_IN_198 WHEN MUX_1024_1_IN_SEL = "0011000110" ELSE
				MUX_1024_1_IN_199 WHEN MUX_1024_1_IN_SEL = "0011000111" ELSE
				MUX_1024_1_IN_200 WHEN MUX_1024_1_IN_SEL = "0011001000" ELSE
				MUX_1024_1_IN_201 WHEN MUX_1024_1_IN_SEL = "0011001001" ELSE
				MUX_1024_1_IN_202 WHEN MUX_1024_1_IN_SEL = "0011001010" ELSE
				MUX_1024_1_IN_203 WHEN MUX_1024_1_IN_SEL = "0011001011" ELSE
				MUX_1024_1_IN_204 WHEN MUX_1024_1_IN_SEL = "0011001100" ELSE
				MUX_1024_1_IN_205 WHEN MUX_1024_1_IN_SEL = "0011001101" ELSE
				MUX_1024_1_IN_206 WHEN MUX_1024_1_IN_SEL = "0011001110" ELSE
				MUX_1024_1_IN_207 WHEN MUX_1024_1_IN_SEL = "0011001111" ELSE
				MUX_1024_1_IN_208 WHEN MUX_1024_1_IN_SEL = "0011010000" ELSE
				MUX_1024_1_IN_209 WHEN MUX_1024_1_IN_SEL = "0011010001" ELSE
				MUX_1024_1_IN_210 WHEN MUX_1024_1_IN_SEL = "0011010010" ELSE
				MUX_1024_1_IN_211 WHEN MUX_1024_1_IN_SEL = "0011010011" ELSE
				MUX_1024_1_IN_212 WHEN MUX_1024_1_IN_SEL = "0011010100" ELSE
				MUX_1024_1_IN_213 WHEN MUX_1024_1_IN_SEL = "0011010101" ELSE
				MUX_1024_1_IN_214 WHEN MUX_1024_1_IN_SEL = "0011010110" ELSE
				MUX_1024_1_IN_215 WHEN MUX_1024_1_IN_SEL = "0011010111" ELSE
				MUX_1024_1_IN_216 WHEN MUX_1024_1_IN_SEL = "0011011000" ELSE
				MUX_1024_1_IN_217 WHEN MUX_1024_1_IN_SEL = "0011011001" ELSE
				MUX_1024_1_IN_218 WHEN MUX_1024_1_IN_SEL = "0011011010" ELSE
				MUX_1024_1_IN_219 WHEN MUX_1024_1_IN_SEL = "0011011011" ELSE
				MUX_1024_1_IN_220 WHEN MUX_1024_1_IN_SEL = "0011011100" ELSE
				MUX_1024_1_IN_221 WHEN MUX_1024_1_IN_SEL = "0011011101" ELSE
				MUX_1024_1_IN_222 WHEN MUX_1024_1_IN_SEL = "0011011110" ELSE
				MUX_1024_1_IN_223 WHEN MUX_1024_1_IN_SEL = "0011011111" ELSE
				MUX_1024_1_IN_224 WHEN MUX_1024_1_IN_SEL = "0011100000" ELSE
				MUX_1024_1_IN_225 WHEN MUX_1024_1_IN_SEL = "0011100001" ELSE
				MUX_1024_1_IN_226 WHEN MUX_1024_1_IN_SEL = "0011100010" ELSE
				MUX_1024_1_IN_227 WHEN MUX_1024_1_IN_SEL = "0011100011" ELSE
				MUX_1024_1_IN_228 WHEN MUX_1024_1_IN_SEL = "0011100100" ELSE
				MUX_1024_1_IN_229 WHEN MUX_1024_1_IN_SEL = "0011100101" ELSE
				MUX_1024_1_IN_230 WHEN MUX_1024_1_IN_SEL = "0011100110" ELSE
				MUX_1024_1_IN_231 WHEN MUX_1024_1_IN_SEL = "0011100111" ELSE
				MUX_1024_1_IN_232 WHEN MUX_1024_1_IN_SEL = "0011101000" ELSE
				MUX_1024_1_IN_233 WHEN MUX_1024_1_IN_SEL = "0011101001" ELSE
				MUX_1024_1_IN_234 WHEN MUX_1024_1_IN_SEL = "0011101010" ELSE
				MUX_1024_1_IN_235 WHEN MUX_1024_1_IN_SEL = "0011101011" ELSE
				MUX_1024_1_IN_236 WHEN MUX_1024_1_IN_SEL = "0011101100" ELSE
				MUX_1024_1_IN_237 WHEN MUX_1024_1_IN_SEL = "0011101101" ELSE
				MUX_1024_1_IN_238 WHEN MUX_1024_1_IN_SEL = "0011101110" ELSE
				MUX_1024_1_IN_239 WHEN MUX_1024_1_IN_SEL = "0011101111" ELSE
				MUX_1024_1_IN_240 WHEN MUX_1024_1_IN_SEL = "0011110000" ELSE
				MUX_1024_1_IN_241 WHEN MUX_1024_1_IN_SEL = "0011110001" ELSE
				MUX_1024_1_IN_242 WHEN MUX_1024_1_IN_SEL = "0011110010" ELSE
				MUX_1024_1_IN_243 WHEN MUX_1024_1_IN_SEL = "0011110011" ELSE
				MUX_1024_1_IN_244 WHEN MUX_1024_1_IN_SEL = "0011110100" ELSE
				MUX_1024_1_IN_245 WHEN MUX_1024_1_IN_SEL = "0011110101" ELSE
				MUX_1024_1_IN_246 WHEN MUX_1024_1_IN_SEL = "0011110110" ELSE
				MUX_1024_1_IN_247 WHEN MUX_1024_1_IN_SEL = "0011110111" ELSE
				MUX_1024_1_IN_248 WHEN MUX_1024_1_IN_SEL = "0011111000" ELSE
				MUX_1024_1_IN_249 WHEN MUX_1024_1_IN_SEL = "0011111001" ELSE
				MUX_1024_1_IN_250 WHEN MUX_1024_1_IN_SEL = "0011111010" ELSE
				MUX_1024_1_IN_251 WHEN MUX_1024_1_IN_SEL = "0011111011" ELSE
				MUX_1024_1_IN_252 WHEN MUX_1024_1_IN_SEL = "0011111100" ELSE
				MUX_1024_1_IN_253 WHEN MUX_1024_1_IN_SEL = "0011111101" ELSE
				MUX_1024_1_IN_254 WHEN MUX_1024_1_IN_SEL = "0011111110" ELSE
				MUX_1024_1_IN_255 WHEN MUX_1024_1_IN_SEL = "0011111111" ELSE
				MUX_1024_1_IN_256 WHEN MUX_1024_1_IN_SEL = "0100000000" ELSE
				MUX_1024_1_IN_257 WHEN MUX_1024_1_IN_SEL = "0100000001" ELSE
				MUX_1024_1_IN_258 WHEN MUX_1024_1_IN_SEL = "0100000010" ELSE
				MUX_1024_1_IN_259 WHEN MUX_1024_1_IN_SEL = "0100000011" ELSE
				MUX_1024_1_IN_260 WHEN MUX_1024_1_IN_SEL = "0100000100" ELSE
				MUX_1024_1_IN_261 WHEN MUX_1024_1_IN_SEL = "0100000101" ELSE
				MUX_1024_1_IN_262 WHEN MUX_1024_1_IN_SEL = "0100000110" ELSE
				MUX_1024_1_IN_263 WHEN MUX_1024_1_IN_SEL = "0100000111" ELSE
				MUX_1024_1_IN_264 WHEN MUX_1024_1_IN_SEL = "0100001000" ELSE
				MUX_1024_1_IN_265 WHEN MUX_1024_1_IN_SEL = "0100001001" ELSE
				MUX_1024_1_IN_266 WHEN MUX_1024_1_IN_SEL = "0100001010" ELSE
				MUX_1024_1_IN_267 WHEN MUX_1024_1_IN_SEL = "0100001011" ELSE
				MUX_1024_1_IN_268 WHEN MUX_1024_1_IN_SEL = "0100001100" ELSE
				MUX_1024_1_IN_269 WHEN MUX_1024_1_IN_SEL = "0100001101" ELSE
				MUX_1024_1_IN_270 WHEN MUX_1024_1_IN_SEL = "0100001110" ELSE
				MUX_1024_1_IN_271 WHEN MUX_1024_1_IN_SEL = "0100001111" ELSE
				MUX_1024_1_IN_272 WHEN MUX_1024_1_IN_SEL = "0100010000" ELSE
				MUX_1024_1_IN_273 WHEN MUX_1024_1_IN_SEL = "0100010001" ELSE
				MUX_1024_1_IN_274 WHEN MUX_1024_1_IN_SEL = "0100010010" ELSE
				MUX_1024_1_IN_275 WHEN MUX_1024_1_IN_SEL = "0100010011" ELSE
				MUX_1024_1_IN_276 WHEN MUX_1024_1_IN_SEL = "0100010100" ELSE
				MUX_1024_1_IN_277 WHEN MUX_1024_1_IN_SEL = "0100010101" ELSE
				MUX_1024_1_IN_278 WHEN MUX_1024_1_IN_SEL = "0100010110" ELSE
				MUX_1024_1_IN_279 WHEN MUX_1024_1_IN_SEL = "0100010111" ELSE
				MUX_1024_1_IN_280 WHEN MUX_1024_1_IN_SEL = "0100011000" ELSE
				MUX_1024_1_IN_281 WHEN MUX_1024_1_IN_SEL = "0100011001" ELSE
				MUX_1024_1_IN_282 WHEN MUX_1024_1_IN_SEL = "0100011010" ELSE
				MUX_1024_1_IN_283 WHEN MUX_1024_1_IN_SEL = "0100011011" ELSE
				MUX_1024_1_IN_284 WHEN MUX_1024_1_IN_SEL = "0100011100" ELSE
				MUX_1024_1_IN_285 WHEN MUX_1024_1_IN_SEL = "0100011101" ELSE
				MUX_1024_1_IN_286 WHEN MUX_1024_1_IN_SEL = "0100011110" ELSE
				MUX_1024_1_IN_287 WHEN MUX_1024_1_IN_SEL = "0100011111" ELSE
				MUX_1024_1_IN_288 WHEN MUX_1024_1_IN_SEL = "0100100000" ELSE
				MUX_1024_1_IN_289 WHEN MUX_1024_1_IN_SEL = "0100100001" ELSE
				MUX_1024_1_IN_290 WHEN MUX_1024_1_IN_SEL = "0100100010" ELSE
				MUX_1024_1_IN_291 WHEN MUX_1024_1_IN_SEL = "0100100011" ELSE
				MUX_1024_1_IN_292 WHEN MUX_1024_1_IN_SEL = "0100100100" ELSE
				MUX_1024_1_IN_293 WHEN MUX_1024_1_IN_SEL = "0100100101" ELSE
				MUX_1024_1_IN_294 WHEN MUX_1024_1_IN_SEL = "0100100110" ELSE
				MUX_1024_1_IN_295 WHEN MUX_1024_1_IN_SEL = "0100100111" ELSE
				MUX_1024_1_IN_296 WHEN MUX_1024_1_IN_SEL = "0100101000" ELSE
				MUX_1024_1_IN_297 WHEN MUX_1024_1_IN_SEL = "0100101001" ELSE
				MUX_1024_1_IN_298 WHEN MUX_1024_1_IN_SEL = "0100101010" ELSE
				MUX_1024_1_IN_299 WHEN MUX_1024_1_IN_SEL = "0100101011" ELSE
				MUX_1024_1_IN_300 WHEN MUX_1024_1_IN_SEL = "0100101100" ELSE
				MUX_1024_1_IN_301 WHEN MUX_1024_1_IN_SEL = "0100101101" ELSE
				MUX_1024_1_IN_302 WHEN MUX_1024_1_IN_SEL = "0100101110" ELSE
				MUX_1024_1_IN_303 WHEN MUX_1024_1_IN_SEL = "0100101111" ELSE
				MUX_1024_1_IN_304 WHEN MUX_1024_1_IN_SEL = "0100110000" ELSE
				MUX_1024_1_IN_305 WHEN MUX_1024_1_IN_SEL = "0100110001" ELSE
				MUX_1024_1_IN_306 WHEN MUX_1024_1_IN_SEL = "0100110010" ELSE
				MUX_1024_1_IN_307 WHEN MUX_1024_1_IN_SEL = "0100110011" ELSE
				MUX_1024_1_IN_308 WHEN MUX_1024_1_IN_SEL = "0100110100" ELSE
				MUX_1024_1_IN_309 WHEN MUX_1024_1_IN_SEL = "0100110101" ELSE
				MUX_1024_1_IN_310 WHEN MUX_1024_1_IN_SEL = "0100110110" ELSE
				MUX_1024_1_IN_311 WHEN MUX_1024_1_IN_SEL = "0100110111" ELSE
				MUX_1024_1_IN_312 WHEN MUX_1024_1_IN_SEL = "0100111000" ELSE
				MUX_1024_1_IN_313 WHEN MUX_1024_1_IN_SEL = "0100111001" ELSE
				MUX_1024_1_IN_314 WHEN MUX_1024_1_IN_SEL = "0100111010" ELSE
				MUX_1024_1_IN_315 WHEN MUX_1024_1_IN_SEL = "0100111011" ELSE
				MUX_1024_1_IN_316 WHEN MUX_1024_1_IN_SEL = "0100111100" ELSE
				MUX_1024_1_IN_317 WHEN MUX_1024_1_IN_SEL = "0100111101" ELSE
				MUX_1024_1_IN_318 WHEN MUX_1024_1_IN_SEL = "0100111110" ELSE
				MUX_1024_1_IN_319 WHEN MUX_1024_1_IN_SEL = "0100111111" ELSE
				MUX_1024_1_IN_320 WHEN MUX_1024_1_IN_SEL = "0101000000" ELSE
				MUX_1024_1_IN_321 WHEN MUX_1024_1_IN_SEL = "0101000001" ELSE
				MUX_1024_1_IN_322 WHEN MUX_1024_1_IN_SEL = "0101000010" ELSE
				MUX_1024_1_IN_323 WHEN MUX_1024_1_IN_SEL = "0101000011" ELSE
				MUX_1024_1_IN_324 WHEN MUX_1024_1_IN_SEL = "0101000100" ELSE
				MUX_1024_1_IN_325 WHEN MUX_1024_1_IN_SEL = "0101000101" ELSE
				MUX_1024_1_IN_326 WHEN MUX_1024_1_IN_SEL = "0101000110" ELSE
				MUX_1024_1_IN_327 WHEN MUX_1024_1_IN_SEL = "0101000111" ELSE
				MUX_1024_1_IN_328 WHEN MUX_1024_1_IN_SEL = "0101001000" ELSE
				MUX_1024_1_IN_329 WHEN MUX_1024_1_IN_SEL = "0101001001" ELSE
				MUX_1024_1_IN_330 WHEN MUX_1024_1_IN_SEL = "0101001010" ELSE
				MUX_1024_1_IN_331 WHEN MUX_1024_1_IN_SEL = "0101001011" ELSE
				MUX_1024_1_IN_332 WHEN MUX_1024_1_IN_SEL = "0101001100" ELSE
				MUX_1024_1_IN_333 WHEN MUX_1024_1_IN_SEL = "0101001101" ELSE
				MUX_1024_1_IN_334 WHEN MUX_1024_1_IN_SEL = "0101001110" ELSE
				MUX_1024_1_IN_335 WHEN MUX_1024_1_IN_SEL = "0101001111" ELSE
				MUX_1024_1_IN_336 WHEN MUX_1024_1_IN_SEL = "0101010000" ELSE
				MUX_1024_1_IN_337 WHEN MUX_1024_1_IN_SEL = "0101010001" ELSE
				MUX_1024_1_IN_338 WHEN MUX_1024_1_IN_SEL = "0101010010" ELSE
				MUX_1024_1_IN_339 WHEN MUX_1024_1_IN_SEL = "0101010011" ELSE
				MUX_1024_1_IN_340 WHEN MUX_1024_1_IN_SEL = "0101010100" ELSE
				MUX_1024_1_IN_341 WHEN MUX_1024_1_IN_SEL = "0101010101" ELSE
				MUX_1024_1_IN_342 WHEN MUX_1024_1_IN_SEL = "0101010110" ELSE
				MUX_1024_1_IN_343 WHEN MUX_1024_1_IN_SEL = "0101010111" ELSE
				MUX_1024_1_IN_344 WHEN MUX_1024_1_IN_SEL = "0101011000" ELSE
				MUX_1024_1_IN_345 WHEN MUX_1024_1_IN_SEL = "0101011001" ELSE
				MUX_1024_1_IN_346 WHEN MUX_1024_1_IN_SEL = "0101011010" ELSE
				MUX_1024_1_IN_347 WHEN MUX_1024_1_IN_SEL = "0101011011" ELSE
				MUX_1024_1_IN_348 WHEN MUX_1024_1_IN_SEL = "0101011100" ELSE
				MUX_1024_1_IN_349 WHEN MUX_1024_1_IN_SEL = "0101011101" ELSE
				MUX_1024_1_IN_350 WHEN MUX_1024_1_IN_SEL = "0101011110" ELSE
				MUX_1024_1_IN_351 WHEN MUX_1024_1_IN_SEL = "0101011111" ELSE
				MUX_1024_1_IN_352 WHEN MUX_1024_1_IN_SEL = "0101100000" ELSE
				MUX_1024_1_IN_353 WHEN MUX_1024_1_IN_SEL = "0101100001" ELSE
				MUX_1024_1_IN_354 WHEN MUX_1024_1_IN_SEL = "0101100010" ELSE
				MUX_1024_1_IN_355 WHEN MUX_1024_1_IN_SEL = "0101100011" ELSE
				MUX_1024_1_IN_356 WHEN MUX_1024_1_IN_SEL = "0101100100" ELSE
				MUX_1024_1_IN_357 WHEN MUX_1024_1_IN_SEL = "0101100101" ELSE
				MUX_1024_1_IN_358 WHEN MUX_1024_1_IN_SEL = "0101100110" ELSE
				MUX_1024_1_IN_359 WHEN MUX_1024_1_IN_SEL = "0101100111" ELSE
				MUX_1024_1_IN_360 WHEN MUX_1024_1_IN_SEL = "0101101000" ELSE
				MUX_1024_1_IN_361 WHEN MUX_1024_1_IN_SEL = "0101101001" ELSE
				MUX_1024_1_IN_362 WHEN MUX_1024_1_IN_SEL = "0101101010" ELSE
				MUX_1024_1_IN_363 WHEN MUX_1024_1_IN_SEL = "0101101011" ELSE
				MUX_1024_1_IN_364 WHEN MUX_1024_1_IN_SEL = "0101101100" ELSE
				MUX_1024_1_IN_365 WHEN MUX_1024_1_IN_SEL = "0101101101" ELSE
				MUX_1024_1_IN_366 WHEN MUX_1024_1_IN_SEL = "0101101110" ELSE
				MUX_1024_1_IN_367 WHEN MUX_1024_1_IN_SEL = "0101101111" ELSE
				MUX_1024_1_IN_368 WHEN MUX_1024_1_IN_SEL = "0101110000" ELSE
				MUX_1024_1_IN_369 WHEN MUX_1024_1_IN_SEL = "0101110001" ELSE
				MUX_1024_1_IN_370 WHEN MUX_1024_1_IN_SEL = "0101110010" ELSE
				MUX_1024_1_IN_371 WHEN MUX_1024_1_IN_SEL = "0101110011" ELSE
				MUX_1024_1_IN_372 WHEN MUX_1024_1_IN_SEL = "0101110100" ELSE
				MUX_1024_1_IN_373 WHEN MUX_1024_1_IN_SEL = "0101110101" ELSE
				MUX_1024_1_IN_374 WHEN MUX_1024_1_IN_SEL = "0101110110" ELSE
				MUX_1024_1_IN_375 WHEN MUX_1024_1_IN_SEL = "0101110111" ELSE
				MUX_1024_1_IN_376 WHEN MUX_1024_1_IN_SEL = "0101111000" ELSE
				MUX_1024_1_IN_377 WHEN MUX_1024_1_IN_SEL = "0101111001" ELSE
				MUX_1024_1_IN_378 WHEN MUX_1024_1_IN_SEL = "0101111010" ELSE
				MUX_1024_1_IN_379 WHEN MUX_1024_1_IN_SEL = "0101111011" ELSE
				MUX_1024_1_IN_380 WHEN MUX_1024_1_IN_SEL = "0101111100" ELSE
				MUX_1024_1_IN_381 WHEN MUX_1024_1_IN_SEL = "0101111101" ELSE
				MUX_1024_1_IN_382 WHEN MUX_1024_1_IN_SEL = "0101111110" ELSE
				MUX_1024_1_IN_383 WHEN MUX_1024_1_IN_SEL = "0101111111" ELSE
				MUX_1024_1_IN_384 WHEN MUX_1024_1_IN_SEL = "0110000000" ELSE
				MUX_1024_1_IN_385 WHEN MUX_1024_1_IN_SEL = "0110000001" ELSE
				MUX_1024_1_IN_386 WHEN MUX_1024_1_IN_SEL = "0110000010" ELSE
				MUX_1024_1_IN_387 WHEN MUX_1024_1_IN_SEL = "0110000011" ELSE
				MUX_1024_1_IN_388 WHEN MUX_1024_1_IN_SEL = "0110000100" ELSE
				MUX_1024_1_IN_389 WHEN MUX_1024_1_IN_SEL = "0110000101" ELSE
				MUX_1024_1_IN_390 WHEN MUX_1024_1_IN_SEL = "0110000110" ELSE
				MUX_1024_1_IN_391 WHEN MUX_1024_1_IN_SEL = "0110000111" ELSE
				MUX_1024_1_IN_392 WHEN MUX_1024_1_IN_SEL = "0110001000" ELSE
				MUX_1024_1_IN_393 WHEN MUX_1024_1_IN_SEL = "0110001001" ELSE
				MUX_1024_1_IN_394 WHEN MUX_1024_1_IN_SEL = "0110001010" ELSE
				MUX_1024_1_IN_395 WHEN MUX_1024_1_IN_SEL = "0110001011" ELSE
				MUX_1024_1_IN_396 WHEN MUX_1024_1_IN_SEL = "0110001100" ELSE
				MUX_1024_1_IN_397 WHEN MUX_1024_1_IN_SEL = "0110001101" ELSE
				MUX_1024_1_IN_398 WHEN MUX_1024_1_IN_SEL = "0110001110" ELSE
				MUX_1024_1_IN_399 WHEN MUX_1024_1_IN_SEL = "0110001111" ELSE
				MUX_1024_1_IN_400 WHEN MUX_1024_1_IN_SEL = "0110010000" ELSE
				MUX_1024_1_IN_401 WHEN MUX_1024_1_IN_SEL = "0110010001" ELSE
				MUX_1024_1_IN_402 WHEN MUX_1024_1_IN_SEL = "0110010010" ELSE
				MUX_1024_1_IN_403 WHEN MUX_1024_1_IN_SEL = "0110010011" ELSE
				MUX_1024_1_IN_404 WHEN MUX_1024_1_IN_SEL = "0110010100" ELSE
				MUX_1024_1_IN_405 WHEN MUX_1024_1_IN_SEL = "0110010101" ELSE
				MUX_1024_1_IN_406 WHEN MUX_1024_1_IN_SEL = "0110010110" ELSE
				MUX_1024_1_IN_407 WHEN MUX_1024_1_IN_SEL = "0110010111" ELSE
				MUX_1024_1_IN_408 WHEN MUX_1024_1_IN_SEL = "0110011000" ELSE
				MUX_1024_1_IN_409 WHEN MUX_1024_1_IN_SEL = "0110011001" ELSE
				MUX_1024_1_IN_410 WHEN MUX_1024_1_IN_SEL = "0110011010" ELSE
				MUX_1024_1_IN_411 WHEN MUX_1024_1_IN_SEL = "0110011011" ELSE
				MUX_1024_1_IN_412 WHEN MUX_1024_1_IN_SEL = "0110011100" ELSE
				MUX_1024_1_IN_413 WHEN MUX_1024_1_IN_SEL = "0110011101" ELSE
				MUX_1024_1_IN_414 WHEN MUX_1024_1_IN_SEL = "0110011110" ELSE
				MUX_1024_1_IN_415 WHEN MUX_1024_1_IN_SEL = "0110011111" ELSE
				MUX_1024_1_IN_416 WHEN MUX_1024_1_IN_SEL = "0110100000" ELSE
				MUX_1024_1_IN_417 WHEN MUX_1024_1_IN_SEL = "0110100001" ELSE
				MUX_1024_1_IN_418 WHEN MUX_1024_1_IN_SEL = "0110100010" ELSE
				MUX_1024_1_IN_419 WHEN MUX_1024_1_IN_SEL = "0110100011" ELSE
				MUX_1024_1_IN_420 WHEN MUX_1024_1_IN_SEL = "0110100100" ELSE
				MUX_1024_1_IN_421 WHEN MUX_1024_1_IN_SEL = "0110100101" ELSE
				MUX_1024_1_IN_422 WHEN MUX_1024_1_IN_SEL = "0110100110" ELSE
				MUX_1024_1_IN_423 WHEN MUX_1024_1_IN_SEL = "0110100111" ELSE
				MUX_1024_1_IN_424 WHEN MUX_1024_1_IN_SEL = "0110101000" ELSE
				MUX_1024_1_IN_425 WHEN MUX_1024_1_IN_SEL = "0110101001" ELSE
				MUX_1024_1_IN_426 WHEN MUX_1024_1_IN_SEL = "0110101010" ELSE
				MUX_1024_1_IN_427 WHEN MUX_1024_1_IN_SEL = "0110101011" ELSE
				MUX_1024_1_IN_428 WHEN MUX_1024_1_IN_SEL = "0110101100" ELSE
				MUX_1024_1_IN_429 WHEN MUX_1024_1_IN_SEL = "0110101101" ELSE
				MUX_1024_1_IN_430 WHEN MUX_1024_1_IN_SEL = "0110101110" ELSE
				MUX_1024_1_IN_431 WHEN MUX_1024_1_IN_SEL = "0110101111" ELSE
				MUX_1024_1_IN_432 WHEN MUX_1024_1_IN_SEL = "0110110000" ELSE
				MUX_1024_1_IN_433 WHEN MUX_1024_1_IN_SEL = "0110110001" ELSE
				MUX_1024_1_IN_434 WHEN MUX_1024_1_IN_SEL = "0110110010" ELSE
				MUX_1024_1_IN_435 WHEN MUX_1024_1_IN_SEL = "0110110011" ELSE
				MUX_1024_1_IN_436 WHEN MUX_1024_1_IN_SEL = "0110110100" ELSE
				MUX_1024_1_IN_437 WHEN MUX_1024_1_IN_SEL = "0110110101" ELSE
				MUX_1024_1_IN_438 WHEN MUX_1024_1_IN_SEL = "0110110110" ELSE
				MUX_1024_1_IN_439 WHEN MUX_1024_1_IN_SEL = "0110110111" ELSE
				MUX_1024_1_IN_440 WHEN MUX_1024_1_IN_SEL = "0110111000" ELSE
				MUX_1024_1_IN_441 WHEN MUX_1024_1_IN_SEL = "0110111001" ELSE
				MUX_1024_1_IN_442 WHEN MUX_1024_1_IN_SEL = "0110111010" ELSE
				MUX_1024_1_IN_443 WHEN MUX_1024_1_IN_SEL = "0110111011" ELSE
				MUX_1024_1_IN_444 WHEN MUX_1024_1_IN_SEL = "0110111100" ELSE
				MUX_1024_1_IN_445 WHEN MUX_1024_1_IN_SEL = "0110111101" ELSE
				MUX_1024_1_IN_446 WHEN MUX_1024_1_IN_SEL = "0110111110" ELSE
				MUX_1024_1_IN_447 WHEN MUX_1024_1_IN_SEL = "0110111111" ELSE
				MUX_1024_1_IN_448 WHEN MUX_1024_1_IN_SEL = "0111000000" ELSE
				MUX_1024_1_IN_449 WHEN MUX_1024_1_IN_SEL = "0111000001" ELSE
				MUX_1024_1_IN_450 WHEN MUX_1024_1_IN_SEL = "0111000010" ELSE
				MUX_1024_1_IN_451 WHEN MUX_1024_1_IN_SEL = "0111000011" ELSE
				MUX_1024_1_IN_452 WHEN MUX_1024_1_IN_SEL = "0111000100" ELSE
				MUX_1024_1_IN_453 WHEN MUX_1024_1_IN_SEL = "0111000101" ELSE
				MUX_1024_1_IN_454 WHEN MUX_1024_1_IN_SEL = "0111000110" ELSE
				MUX_1024_1_IN_455 WHEN MUX_1024_1_IN_SEL = "0111000111" ELSE
				MUX_1024_1_IN_456 WHEN MUX_1024_1_IN_SEL = "0111001000" ELSE
				MUX_1024_1_IN_457 WHEN MUX_1024_1_IN_SEL = "0111001001" ELSE
				MUX_1024_1_IN_458 WHEN MUX_1024_1_IN_SEL = "0111001010" ELSE
				MUX_1024_1_IN_459 WHEN MUX_1024_1_IN_SEL = "0111001011" ELSE
				MUX_1024_1_IN_460 WHEN MUX_1024_1_IN_SEL = "0111001100" ELSE
				MUX_1024_1_IN_461 WHEN MUX_1024_1_IN_SEL = "0111001101" ELSE
				MUX_1024_1_IN_462 WHEN MUX_1024_1_IN_SEL = "0111001110" ELSE
				MUX_1024_1_IN_463 WHEN MUX_1024_1_IN_SEL = "0111001111" ELSE
				MUX_1024_1_IN_464 WHEN MUX_1024_1_IN_SEL = "0111010000" ELSE
				MUX_1024_1_IN_465 WHEN MUX_1024_1_IN_SEL = "0111010001" ELSE
				MUX_1024_1_IN_466 WHEN MUX_1024_1_IN_SEL = "0111010010" ELSE
				MUX_1024_1_IN_467 WHEN MUX_1024_1_IN_SEL = "0111010011" ELSE
				MUX_1024_1_IN_468 WHEN MUX_1024_1_IN_SEL = "0111010100" ELSE
				MUX_1024_1_IN_469 WHEN MUX_1024_1_IN_SEL = "0111010101" ELSE
				MUX_1024_1_IN_470 WHEN MUX_1024_1_IN_SEL = "0111010110" ELSE
				MUX_1024_1_IN_471 WHEN MUX_1024_1_IN_SEL = "0111010111" ELSE
				MUX_1024_1_IN_472 WHEN MUX_1024_1_IN_SEL = "0111011000" ELSE
				MUX_1024_1_IN_473 WHEN MUX_1024_1_IN_SEL = "0111011001" ELSE
				MUX_1024_1_IN_474 WHEN MUX_1024_1_IN_SEL = "0111011010" ELSE
				MUX_1024_1_IN_475 WHEN MUX_1024_1_IN_SEL = "0111011011" ELSE
				MUX_1024_1_IN_476 WHEN MUX_1024_1_IN_SEL = "0111011100" ELSE
				MUX_1024_1_IN_477 WHEN MUX_1024_1_IN_SEL = "0111011101" ELSE
				MUX_1024_1_IN_478 WHEN MUX_1024_1_IN_SEL = "0111011110" ELSE
				MUX_1024_1_IN_479 WHEN MUX_1024_1_IN_SEL = "0111011111" ELSE
				MUX_1024_1_IN_480 WHEN MUX_1024_1_IN_SEL = "0111100000" ELSE
				MUX_1024_1_IN_481 WHEN MUX_1024_1_IN_SEL = "0111100001" ELSE
				MUX_1024_1_IN_482 WHEN MUX_1024_1_IN_SEL = "0111100010" ELSE
				MUX_1024_1_IN_483 WHEN MUX_1024_1_IN_SEL = "0111100011" ELSE
				MUX_1024_1_IN_484 WHEN MUX_1024_1_IN_SEL = "0111100100" ELSE
				MUX_1024_1_IN_485 WHEN MUX_1024_1_IN_SEL = "0111100101" ELSE
				MUX_1024_1_IN_486 WHEN MUX_1024_1_IN_SEL = "0111100110" ELSE
				MUX_1024_1_IN_487 WHEN MUX_1024_1_IN_SEL = "0111100111" ELSE
				MUX_1024_1_IN_488 WHEN MUX_1024_1_IN_SEL = "0111101000" ELSE
				MUX_1024_1_IN_489 WHEN MUX_1024_1_IN_SEL = "0111101001" ELSE
				MUX_1024_1_IN_490 WHEN MUX_1024_1_IN_SEL = "0111101010" ELSE
				MUX_1024_1_IN_491 WHEN MUX_1024_1_IN_SEL = "0111101011" ELSE
				MUX_1024_1_IN_492 WHEN MUX_1024_1_IN_SEL = "0111101100" ELSE
				MUX_1024_1_IN_493 WHEN MUX_1024_1_IN_SEL = "0111101101" ELSE
				MUX_1024_1_IN_494 WHEN MUX_1024_1_IN_SEL = "0111101110" ELSE
				MUX_1024_1_IN_495 WHEN MUX_1024_1_IN_SEL = "0111101111" ELSE
				MUX_1024_1_IN_496 WHEN MUX_1024_1_IN_SEL = "0111110000" ELSE
				MUX_1024_1_IN_497 WHEN MUX_1024_1_IN_SEL = "0111110001" ELSE
				MUX_1024_1_IN_498 WHEN MUX_1024_1_IN_SEL = "0111110010" ELSE
				MUX_1024_1_IN_499 WHEN MUX_1024_1_IN_SEL = "0111110011" ELSE
				MUX_1024_1_IN_500 WHEN MUX_1024_1_IN_SEL = "0111110100" ELSE
				MUX_1024_1_IN_501 WHEN MUX_1024_1_IN_SEL = "0111110101" ELSE
				MUX_1024_1_IN_502 WHEN MUX_1024_1_IN_SEL = "0111110110" ELSE
				MUX_1024_1_IN_503 WHEN MUX_1024_1_IN_SEL = "0111110111" ELSE
				MUX_1024_1_IN_504 WHEN MUX_1024_1_IN_SEL = "0111111000" ELSE
				MUX_1024_1_IN_505 WHEN MUX_1024_1_IN_SEL = "0111111001" ELSE
				MUX_1024_1_IN_506 WHEN MUX_1024_1_IN_SEL = "0111111010" ELSE
				MUX_1024_1_IN_507 WHEN MUX_1024_1_IN_SEL = "0111111011" ELSE
				MUX_1024_1_IN_508 WHEN MUX_1024_1_IN_SEL = "0111111100" ELSE
				MUX_1024_1_IN_509 WHEN MUX_1024_1_IN_SEL = "0111111101" ELSE
				MUX_1024_1_IN_510 WHEN MUX_1024_1_IN_SEL = "0111111110" ELSE
				MUX_1024_1_IN_511 WHEN MUX_1024_1_IN_SEL = "0111111111" ELSE
				MUX_1024_1_IN_512 WHEN MUX_1024_1_IN_SEL = "1000000000" ELSE
				MUX_1024_1_IN_513 WHEN MUX_1024_1_IN_SEL = "1000000001" ELSE
				MUX_1024_1_IN_514 WHEN MUX_1024_1_IN_SEL = "1000000010" ELSE
				MUX_1024_1_IN_515 WHEN MUX_1024_1_IN_SEL = "1000000011" ELSE
				MUX_1024_1_IN_516 WHEN MUX_1024_1_IN_SEL = "1000000100" ELSE
				MUX_1024_1_IN_517 WHEN MUX_1024_1_IN_SEL = "1000000101" ELSE
				MUX_1024_1_IN_518 WHEN MUX_1024_1_IN_SEL = "1000000110" ELSE
				MUX_1024_1_IN_519 WHEN MUX_1024_1_IN_SEL = "1000000111" ELSE
				MUX_1024_1_IN_520 WHEN MUX_1024_1_IN_SEL = "1000001000" ELSE
				MUX_1024_1_IN_521 WHEN MUX_1024_1_IN_SEL = "1000001001" ELSE
				MUX_1024_1_IN_522 WHEN MUX_1024_1_IN_SEL = "1000001010" ELSE
				MUX_1024_1_IN_523 WHEN MUX_1024_1_IN_SEL = "1000001011" ELSE
				MUX_1024_1_IN_524 WHEN MUX_1024_1_IN_SEL = "1000001100" ELSE
				MUX_1024_1_IN_525 WHEN MUX_1024_1_IN_SEL = "1000001101" ELSE
				MUX_1024_1_IN_526 WHEN MUX_1024_1_IN_SEL = "1000001110" ELSE
				MUX_1024_1_IN_527 WHEN MUX_1024_1_IN_SEL = "1000001111" ELSE
				MUX_1024_1_IN_528 WHEN MUX_1024_1_IN_SEL = "1000010000" ELSE
				MUX_1024_1_IN_529 WHEN MUX_1024_1_IN_SEL = "1000010001" ELSE
				MUX_1024_1_IN_530 WHEN MUX_1024_1_IN_SEL = "1000010010" ELSE
				MUX_1024_1_IN_531 WHEN MUX_1024_1_IN_SEL = "1000010011" ELSE
				MUX_1024_1_IN_532 WHEN MUX_1024_1_IN_SEL = "1000010100" ELSE
				MUX_1024_1_IN_533 WHEN MUX_1024_1_IN_SEL = "1000010101" ELSE
				MUX_1024_1_IN_534 WHEN MUX_1024_1_IN_SEL = "1000010110" ELSE
				MUX_1024_1_IN_535 WHEN MUX_1024_1_IN_SEL = "1000010111" ELSE
				MUX_1024_1_IN_536 WHEN MUX_1024_1_IN_SEL = "1000011000" ELSE
				MUX_1024_1_IN_537 WHEN MUX_1024_1_IN_SEL = "1000011001" ELSE
				MUX_1024_1_IN_538 WHEN MUX_1024_1_IN_SEL = "1000011010" ELSE
				MUX_1024_1_IN_539 WHEN MUX_1024_1_IN_SEL = "1000011011" ELSE
				MUX_1024_1_IN_540 WHEN MUX_1024_1_IN_SEL = "1000011100" ELSE
				MUX_1024_1_IN_541 WHEN MUX_1024_1_IN_SEL = "1000011101" ELSE
				MUX_1024_1_IN_542 WHEN MUX_1024_1_IN_SEL = "1000011110" ELSE
				MUX_1024_1_IN_543 WHEN MUX_1024_1_IN_SEL = "1000011111" ELSE
				MUX_1024_1_IN_544 WHEN MUX_1024_1_IN_SEL = "1000100000" ELSE
				MUX_1024_1_IN_545 WHEN MUX_1024_1_IN_SEL = "1000100001" ELSE
				MUX_1024_1_IN_546 WHEN MUX_1024_1_IN_SEL = "1000100010" ELSE
				MUX_1024_1_IN_547 WHEN MUX_1024_1_IN_SEL = "1000100011" ELSE
				MUX_1024_1_IN_548 WHEN MUX_1024_1_IN_SEL = "1000100100" ELSE
				MUX_1024_1_IN_549 WHEN MUX_1024_1_IN_SEL = "1000100101" ELSE
				MUX_1024_1_IN_550 WHEN MUX_1024_1_IN_SEL = "1000100110" ELSE
				MUX_1024_1_IN_551 WHEN MUX_1024_1_IN_SEL = "1000100111" ELSE
				MUX_1024_1_IN_552 WHEN MUX_1024_1_IN_SEL = "1000101000" ELSE
				MUX_1024_1_IN_553 WHEN MUX_1024_1_IN_SEL = "1000101001" ELSE
				MUX_1024_1_IN_554 WHEN MUX_1024_1_IN_SEL = "1000101010" ELSE
				MUX_1024_1_IN_555 WHEN MUX_1024_1_IN_SEL = "1000101011" ELSE
				MUX_1024_1_IN_556 WHEN MUX_1024_1_IN_SEL = "1000101100" ELSE
				MUX_1024_1_IN_557 WHEN MUX_1024_1_IN_SEL = "1000101101" ELSE
				MUX_1024_1_IN_558 WHEN MUX_1024_1_IN_SEL = "1000101110" ELSE
				MUX_1024_1_IN_559 WHEN MUX_1024_1_IN_SEL = "1000101111" ELSE
				MUX_1024_1_IN_560 WHEN MUX_1024_1_IN_SEL = "1000110000" ELSE
				MUX_1024_1_IN_561 WHEN MUX_1024_1_IN_SEL = "1000110001" ELSE
				MUX_1024_1_IN_562 WHEN MUX_1024_1_IN_SEL = "1000110010" ELSE
				MUX_1024_1_IN_563 WHEN MUX_1024_1_IN_SEL = "1000110011" ELSE
				MUX_1024_1_IN_564 WHEN MUX_1024_1_IN_SEL = "1000110100" ELSE
				MUX_1024_1_IN_565 WHEN MUX_1024_1_IN_SEL = "1000110101" ELSE
				MUX_1024_1_IN_566 WHEN MUX_1024_1_IN_SEL = "1000110110" ELSE
				MUX_1024_1_IN_567 WHEN MUX_1024_1_IN_SEL = "1000110111" ELSE
				MUX_1024_1_IN_568 WHEN MUX_1024_1_IN_SEL = "1000111000" ELSE
				MUX_1024_1_IN_569 WHEN MUX_1024_1_IN_SEL = "1000111001" ELSE
				MUX_1024_1_IN_570 WHEN MUX_1024_1_IN_SEL = "1000111010" ELSE
				MUX_1024_1_IN_571 WHEN MUX_1024_1_IN_SEL = "1000111011" ELSE
				MUX_1024_1_IN_572 WHEN MUX_1024_1_IN_SEL = "1000111100" ELSE
				MUX_1024_1_IN_573 WHEN MUX_1024_1_IN_SEL = "1000111101" ELSE
				MUX_1024_1_IN_574 WHEN MUX_1024_1_IN_SEL = "1000111110" ELSE
				MUX_1024_1_IN_575 WHEN MUX_1024_1_IN_SEL = "1000111111" ELSE
				MUX_1024_1_IN_576 WHEN MUX_1024_1_IN_SEL = "1001000000" ELSE
				MUX_1024_1_IN_577 WHEN MUX_1024_1_IN_SEL = "1001000001" ELSE
				MUX_1024_1_IN_578 WHEN MUX_1024_1_IN_SEL = "1001000010" ELSE
				MUX_1024_1_IN_579 WHEN MUX_1024_1_IN_SEL = "1001000011" ELSE
				MUX_1024_1_IN_580 WHEN MUX_1024_1_IN_SEL = "1001000100" ELSE
				MUX_1024_1_IN_581 WHEN MUX_1024_1_IN_SEL = "1001000101" ELSE
				MUX_1024_1_IN_582 WHEN MUX_1024_1_IN_SEL = "1001000110" ELSE
				MUX_1024_1_IN_583 WHEN MUX_1024_1_IN_SEL = "1001000111" ELSE
				MUX_1024_1_IN_584 WHEN MUX_1024_1_IN_SEL = "1001001000" ELSE
				MUX_1024_1_IN_585 WHEN MUX_1024_1_IN_SEL = "1001001001" ELSE
				MUX_1024_1_IN_586 WHEN MUX_1024_1_IN_SEL = "1001001010" ELSE
				MUX_1024_1_IN_587 WHEN MUX_1024_1_IN_SEL = "1001001011" ELSE
				MUX_1024_1_IN_588 WHEN MUX_1024_1_IN_SEL = "1001001100" ELSE
				MUX_1024_1_IN_589 WHEN MUX_1024_1_IN_SEL = "1001001101" ELSE
				MUX_1024_1_IN_590 WHEN MUX_1024_1_IN_SEL = "1001001110" ELSE
				MUX_1024_1_IN_591 WHEN MUX_1024_1_IN_SEL = "1001001111" ELSE
				MUX_1024_1_IN_592 WHEN MUX_1024_1_IN_SEL = "1001010000" ELSE
				MUX_1024_1_IN_593 WHEN MUX_1024_1_IN_SEL = "1001010001" ELSE
				MUX_1024_1_IN_594 WHEN MUX_1024_1_IN_SEL = "1001010010" ELSE
				MUX_1024_1_IN_595 WHEN MUX_1024_1_IN_SEL = "1001010011" ELSE
				MUX_1024_1_IN_596 WHEN MUX_1024_1_IN_SEL = "1001010100" ELSE
				MUX_1024_1_IN_597 WHEN MUX_1024_1_IN_SEL = "1001010101" ELSE
				MUX_1024_1_IN_598 WHEN MUX_1024_1_IN_SEL = "1001010110" ELSE
				MUX_1024_1_IN_599 WHEN MUX_1024_1_IN_SEL = "1001010111" ELSE
				MUX_1024_1_IN_600 WHEN MUX_1024_1_IN_SEL = "1001011000" ELSE
				MUX_1024_1_IN_601 WHEN MUX_1024_1_IN_SEL = "1001011001" ELSE
				MUX_1024_1_IN_602 WHEN MUX_1024_1_IN_SEL = "1001011010" ELSE
				MUX_1024_1_IN_603 WHEN MUX_1024_1_IN_SEL = "1001011011" ELSE
				MUX_1024_1_IN_604 WHEN MUX_1024_1_IN_SEL = "1001011100" ELSE
				MUX_1024_1_IN_605 WHEN MUX_1024_1_IN_SEL = "1001011101" ELSE
				MUX_1024_1_IN_606 WHEN MUX_1024_1_IN_SEL = "1001011110" ELSE
				MUX_1024_1_IN_607 WHEN MUX_1024_1_IN_SEL = "1001011111" ELSE
				MUX_1024_1_IN_608 WHEN MUX_1024_1_IN_SEL = "1001100000" ELSE
				MUX_1024_1_IN_609 WHEN MUX_1024_1_IN_SEL = "1001100001" ELSE
				MUX_1024_1_IN_610 WHEN MUX_1024_1_IN_SEL = "1001100010" ELSE
				MUX_1024_1_IN_611 WHEN MUX_1024_1_IN_SEL = "1001100011" ELSE
				MUX_1024_1_IN_612 WHEN MUX_1024_1_IN_SEL = "1001100100" ELSE
				MUX_1024_1_IN_613 WHEN MUX_1024_1_IN_SEL = "1001100101" ELSE
				MUX_1024_1_IN_614 WHEN MUX_1024_1_IN_SEL = "1001100110" ELSE
				MUX_1024_1_IN_615 WHEN MUX_1024_1_IN_SEL = "1001100111" ELSE
				MUX_1024_1_IN_616 WHEN MUX_1024_1_IN_SEL = "1001101000" ELSE
				MUX_1024_1_IN_617 WHEN MUX_1024_1_IN_SEL = "1001101001" ELSE
				MUX_1024_1_IN_618 WHEN MUX_1024_1_IN_SEL = "1001101010" ELSE
				MUX_1024_1_IN_619 WHEN MUX_1024_1_IN_SEL = "1001101011" ELSE
				MUX_1024_1_IN_620 WHEN MUX_1024_1_IN_SEL = "1001101100" ELSE
				MUX_1024_1_IN_621 WHEN MUX_1024_1_IN_SEL = "1001101101" ELSE
				MUX_1024_1_IN_622 WHEN MUX_1024_1_IN_SEL = "1001101110" ELSE
				MUX_1024_1_IN_623 WHEN MUX_1024_1_IN_SEL = "1001101111" ELSE
				MUX_1024_1_IN_624 WHEN MUX_1024_1_IN_SEL = "1001110000" ELSE
				MUX_1024_1_IN_625 WHEN MUX_1024_1_IN_SEL = "1001110001" ELSE
				MUX_1024_1_IN_626 WHEN MUX_1024_1_IN_SEL = "1001110010" ELSE
				MUX_1024_1_IN_627 WHEN MUX_1024_1_IN_SEL = "1001110011" ELSE
				MUX_1024_1_IN_628 WHEN MUX_1024_1_IN_SEL = "1001110100" ELSE
				MUX_1024_1_IN_629 WHEN MUX_1024_1_IN_SEL = "1001110101" ELSE
				MUX_1024_1_IN_630 WHEN MUX_1024_1_IN_SEL = "1001110110" ELSE
				MUX_1024_1_IN_631 WHEN MUX_1024_1_IN_SEL = "1001110111" ELSE
				MUX_1024_1_IN_632 WHEN MUX_1024_1_IN_SEL = "1001111000" ELSE
				MUX_1024_1_IN_633 WHEN MUX_1024_1_IN_SEL = "1001111001" ELSE
				MUX_1024_1_IN_634 WHEN MUX_1024_1_IN_SEL = "1001111010" ELSE
				MUX_1024_1_IN_635 WHEN MUX_1024_1_IN_SEL = "1001111011" ELSE
				MUX_1024_1_IN_636 WHEN MUX_1024_1_IN_SEL = "1001111100" ELSE
				MUX_1024_1_IN_637 WHEN MUX_1024_1_IN_SEL = "1001111101" ELSE
				MUX_1024_1_IN_638 WHEN MUX_1024_1_IN_SEL = "1001111110" ELSE
				MUX_1024_1_IN_639 WHEN MUX_1024_1_IN_SEL = "1001111111" ELSE
				MUX_1024_1_IN_640 WHEN MUX_1024_1_IN_SEL = "1010000000" ELSE
				MUX_1024_1_IN_641 WHEN MUX_1024_1_IN_SEL = "1010000001" ELSE
				MUX_1024_1_IN_642 WHEN MUX_1024_1_IN_SEL = "1010000010" ELSE
				MUX_1024_1_IN_643 WHEN MUX_1024_1_IN_SEL = "1010000011" ELSE
				MUX_1024_1_IN_644 WHEN MUX_1024_1_IN_SEL = "1010000100" ELSE
				MUX_1024_1_IN_645 WHEN MUX_1024_1_IN_SEL = "1010000101" ELSE
				MUX_1024_1_IN_646 WHEN MUX_1024_1_IN_SEL = "1010000110" ELSE
				MUX_1024_1_IN_647 WHEN MUX_1024_1_IN_SEL = "1010000111" ELSE
				MUX_1024_1_IN_648 WHEN MUX_1024_1_IN_SEL = "1010001000" ELSE
				MUX_1024_1_IN_649 WHEN MUX_1024_1_IN_SEL = "1010001001" ELSE
				MUX_1024_1_IN_650 WHEN MUX_1024_1_IN_SEL = "1010001010" ELSE
				MUX_1024_1_IN_651 WHEN MUX_1024_1_IN_SEL = "1010001011" ELSE
				MUX_1024_1_IN_652 WHEN MUX_1024_1_IN_SEL = "1010001100" ELSE
				MUX_1024_1_IN_653 WHEN MUX_1024_1_IN_SEL = "1010001101" ELSE
				MUX_1024_1_IN_654 WHEN MUX_1024_1_IN_SEL = "1010001110" ELSE
				MUX_1024_1_IN_655 WHEN MUX_1024_1_IN_SEL = "1010001111" ELSE
				MUX_1024_1_IN_656 WHEN MUX_1024_1_IN_SEL = "1010010000" ELSE
				MUX_1024_1_IN_657 WHEN MUX_1024_1_IN_SEL = "1010010001" ELSE
				MUX_1024_1_IN_658 WHEN MUX_1024_1_IN_SEL = "1010010010" ELSE
				MUX_1024_1_IN_659 WHEN MUX_1024_1_IN_SEL = "1010010011" ELSE
				MUX_1024_1_IN_660 WHEN MUX_1024_1_IN_SEL = "1010010100" ELSE
				MUX_1024_1_IN_661 WHEN MUX_1024_1_IN_SEL = "1010010101" ELSE
				MUX_1024_1_IN_662 WHEN MUX_1024_1_IN_SEL = "1010010110" ELSE
				MUX_1024_1_IN_663 WHEN MUX_1024_1_IN_SEL = "1010010111" ELSE
				MUX_1024_1_IN_664 WHEN MUX_1024_1_IN_SEL = "1010011000" ELSE
				MUX_1024_1_IN_665 WHEN MUX_1024_1_IN_SEL = "1010011001" ELSE
				MUX_1024_1_IN_666 WHEN MUX_1024_1_IN_SEL = "1010011010" ELSE
				MUX_1024_1_IN_667 WHEN MUX_1024_1_IN_SEL = "1010011011" ELSE
				MUX_1024_1_IN_668 WHEN MUX_1024_1_IN_SEL = "1010011100" ELSE
				MUX_1024_1_IN_669 WHEN MUX_1024_1_IN_SEL = "1010011101" ELSE
				MUX_1024_1_IN_670 WHEN MUX_1024_1_IN_SEL = "1010011110" ELSE
				MUX_1024_1_IN_671 WHEN MUX_1024_1_IN_SEL = "1010011111" ELSE
				MUX_1024_1_IN_672 WHEN MUX_1024_1_IN_SEL = "1010100000" ELSE
				MUX_1024_1_IN_673 WHEN MUX_1024_1_IN_SEL = "1010100001" ELSE
				MUX_1024_1_IN_674 WHEN MUX_1024_1_IN_SEL = "1010100010" ELSE
				MUX_1024_1_IN_675 WHEN MUX_1024_1_IN_SEL = "1010100011" ELSE
				MUX_1024_1_IN_676 WHEN MUX_1024_1_IN_SEL = "1010100100" ELSE
				MUX_1024_1_IN_677 WHEN MUX_1024_1_IN_SEL = "1010100101" ELSE
				MUX_1024_1_IN_678 WHEN MUX_1024_1_IN_SEL = "1010100110" ELSE
				MUX_1024_1_IN_679 WHEN MUX_1024_1_IN_SEL = "1010100111" ELSE
				MUX_1024_1_IN_680 WHEN MUX_1024_1_IN_SEL = "1010101000" ELSE
				MUX_1024_1_IN_681 WHEN MUX_1024_1_IN_SEL = "1010101001" ELSE
				MUX_1024_1_IN_682 WHEN MUX_1024_1_IN_SEL = "1010101010" ELSE
				MUX_1024_1_IN_683 WHEN MUX_1024_1_IN_SEL = "1010101011" ELSE
				MUX_1024_1_IN_684 WHEN MUX_1024_1_IN_SEL = "1010101100" ELSE
				MUX_1024_1_IN_685 WHEN MUX_1024_1_IN_SEL = "1010101101" ELSE
				MUX_1024_1_IN_686 WHEN MUX_1024_1_IN_SEL = "1010101110" ELSE
				MUX_1024_1_IN_687 WHEN MUX_1024_1_IN_SEL = "1010101111" ELSE
				MUX_1024_1_IN_688 WHEN MUX_1024_1_IN_SEL = "1010110000" ELSE
				MUX_1024_1_IN_689 WHEN MUX_1024_1_IN_SEL = "1010110001" ELSE
				MUX_1024_1_IN_690 WHEN MUX_1024_1_IN_SEL = "1010110010" ELSE
				MUX_1024_1_IN_691 WHEN MUX_1024_1_IN_SEL = "1010110011" ELSE
				MUX_1024_1_IN_692 WHEN MUX_1024_1_IN_SEL = "1010110100" ELSE
				MUX_1024_1_IN_693 WHEN MUX_1024_1_IN_SEL = "1010110101" ELSE
				MUX_1024_1_IN_694 WHEN MUX_1024_1_IN_SEL = "1010110110" ELSE
				MUX_1024_1_IN_695 WHEN MUX_1024_1_IN_SEL = "1010110111" ELSE
				MUX_1024_1_IN_696 WHEN MUX_1024_1_IN_SEL = "1010111000" ELSE
				MUX_1024_1_IN_697 WHEN MUX_1024_1_IN_SEL = "1010111001" ELSE
				MUX_1024_1_IN_698 WHEN MUX_1024_1_IN_SEL = "1010111010" ELSE
				MUX_1024_1_IN_699 WHEN MUX_1024_1_IN_SEL = "1010111011" ELSE
				MUX_1024_1_IN_700 WHEN MUX_1024_1_IN_SEL = "1010111100" ELSE
				MUX_1024_1_IN_701 WHEN MUX_1024_1_IN_SEL = "1010111101" ELSE
				MUX_1024_1_IN_702 WHEN MUX_1024_1_IN_SEL = "1010111110" ELSE
				MUX_1024_1_IN_703 WHEN MUX_1024_1_IN_SEL = "1010111111" ELSE
				MUX_1024_1_IN_704 WHEN MUX_1024_1_IN_SEL = "1011000000" ELSE
				MUX_1024_1_IN_705 WHEN MUX_1024_1_IN_SEL = "1011000001" ELSE
				MUX_1024_1_IN_706 WHEN MUX_1024_1_IN_SEL = "1011000010" ELSE
				MUX_1024_1_IN_707 WHEN MUX_1024_1_IN_SEL = "1011000011" ELSE
				MUX_1024_1_IN_708 WHEN MUX_1024_1_IN_SEL = "1011000100" ELSE
				MUX_1024_1_IN_709 WHEN MUX_1024_1_IN_SEL = "1011000101" ELSE
				MUX_1024_1_IN_710 WHEN MUX_1024_1_IN_SEL = "1011000110" ELSE
				MUX_1024_1_IN_711 WHEN MUX_1024_1_IN_SEL = "1011000111" ELSE
				MUX_1024_1_IN_712 WHEN MUX_1024_1_IN_SEL = "1011001000" ELSE
				MUX_1024_1_IN_713 WHEN MUX_1024_1_IN_SEL = "1011001001" ELSE
				MUX_1024_1_IN_714 WHEN MUX_1024_1_IN_SEL = "1011001010" ELSE
				MUX_1024_1_IN_715 WHEN MUX_1024_1_IN_SEL = "1011001011" ELSE
				MUX_1024_1_IN_716 WHEN MUX_1024_1_IN_SEL = "1011001100" ELSE
				MUX_1024_1_IN_717 WHEN MUX_1024_1_IN_SEL = "1011001101" ELSE
				MUX_1024_1_IN_718 WHEN MUX_1024_1_IN_SEL = "1011001110" ELSE
				MUX_1024_1_IN_719 WHEN MUX_1024_1_IN_SEL = "1011001111" ELSE
				MUX_1024_1_IN_720 WHEN MUX_1024_1_IN_SEL = "1011010000" ELSE
				MUX_1024_1_IN_721 WHEN MUX_1024_1_IN_SEL = "1011010001" ELSE
				MUX_1024_1_IN_722 WHEN MUX_1024_1_IN_SEL = "1011010010" ELSE
				MUX_1024_1_IN_723 WHEN MUX_1024_1_IN_SEL = "1011010011" ELSE
				MUX_1024_1_IN_724 WHEN MUX_1024_1_IN_SEL = "1011010100" ELSE
				MUX_1024_1_IN_725 WHEN MUX_1024_1_IN_SEL = "1011010101" ELSE
				MUX_1024_1_IN_726 WHEN MUX_1024_1_IN_SEL = "1011010110" ELSE
				MUX_1024_1_IN_727 WHEN MUX_1024_1_IN_SEL = "1011010111" ELSE
				MUX_1024_1_IN_728 WHEN MUX_1024_1_IN_SEL = "1011011000" ELSE
				MUX_1024_1_IN_729 WHEN MUX_1024_1_IN_SEL = "1011011001" ELSE
				MUX_1024_1_IN_730 WHEN MUX_1024_1_IN_SEL = "1011011010" ELSE
				MUX_1024_1_IN_731 WHEN MUX_1024_1_IN_SEL = "1011011011" ELSE
				MUX_1024_1_IN_732 WHEN MUX_1024_1_IN_SEL = "1011011100" ELSE
				MUX_1024_1_IN_733 WHEN MUX_1024_1_IN_SEL = "1011011101" ELSE
				MUX_1024_1_IN_734 WHEN MUX_1024_1_IN_SEL = "1011011110" ELSE
				MUX_1024_1_IN_735 WHEN MUX_1024_1_IN_SEL = "1011011111" ELSE
				MUX_1024_1_IN_736 WHEN MUX_1024_1_IN_SEL = "1011100000" ELSE
				MUX_1024_1_IN_737 WHEN MUX_1024_1_IN_SEL = "1011100001" ELSE
				MUX_1024_1_IN_738 WHEN MUX_1024_1_IN_SEL = "1011100010" ELSE
				MUX_1024_1_IN_739 WHEN MUX_1024_1_IN_SEL = "1011100011" ELSE
				MUX_1024_1_IN_740 WHEN MUX_1024_1_IN_SEL = "1011100100" ELSE
				MUX_1024_1_IN_741 WHEN MUX_1024_1_IN_SEL = "1011100101" ELSE
				MUX_1024_1_IN_742 WHEN MUX_1024_1_IN_SEL = "1011100110" ELSE
				MUX_1024_1_IN_743 WHEN MUX_1024_1_IN_SEL = "1011100111" ELSE
				MUX_1024_1_IN_744 WHEN MUX_1024_1_IN_SEL = "1011101000" ELSE
				MUX_1024_1_IN_745 WHEN MUX_1024_1_IN_SEL = "1011101001" ELSE
				MUX_1024_1_IN_746 WHEN MUX_1024_1_IN_SEL = "1011101010" ELSE
				MUX_1024_1_IN_747 WHEN MUX_1024_1_IN_SEL = "1011101011" ELSE
				MUX_1024_1_IN_748 WHEN MUX_1024_1_IN_SEL = "1011101100" ELSE
				MUX_1024_1_IN_749 WHEN MUX_1024_1_IN_SEL = "1011101101" ELSE
				MUX_1024_1_IN_750 WHEN MUX_1024_1_IN_SEL = "1011101110" ELSE
				MUX_1024_1_IN_751 WHEN MUX_1024_1_IN_SEL = "1011101111" ELSE
				MUX_1024_1_IN_752 WHEN MUX_1024_1_IN_SEL = "1011110000" ELSE
				MUX_1024_1_IN_753 WHEN MUX_1024_1_IN_SEL = "1011110001" ELSE
				MUX_1024_1_IN_754 WHEN MUX_1024_1_IN_SEL = "1011110010" ELSE
				MUX_1024_1_IN_755 WHEN MUX_1024_1_IN_SEL = "1011110011" ELSE
				MUX_1024_1_IN_756 WHEN MUX_1024_1_IN_SEL = "1011110100" ELSE
				MUX_1024_1_IN_757 WHEN MUX_1024_1_IN_SEL = "1011110101" ELSE
				MUX_1024_1_IN_758 WHEN MUX_1024_1_IN_SEL = "1011110110" ELSE
				MUX_1024_1_IN_759 WHEN MUX_1024_1_IN_SEL = "1011110111" ELSE
				MUX_1024_1_IN_760 WHEN MUX_1024_1_IN_SEL = "1011111000" ELSE
				MUX_1024_1_IN_761 WHEN MUX_1024_1_IN_SEL = "1011111001" ELSE
				MUX_1024_1_IN_762 WHEN MUX_1024_1_IN_SEL = "1011111010" ELSE
				MUX_1024_1_IN_763 WHEN MUX_1024_1_IN_SEL = "1011111011" ELSE
				MUX_1024_1_IN_764 WHEN MUX_1024_1_IN_SEL = "1011111100" ELSE
				MUX_1024_1_IN_765 WHEN MUX_1024_1_IN_SEL = "1011111101" ELSE
				MUX_1024_1_IN_766 WHEN MUX_1024_1_IN_SEL = "1011111110" ELSE
				MUX_1024_1_IN_767 WHEN MUX_1024_1_IN_SEL = "1011111111" ELSE
				MUX_1024_1_IN_768 WHEN MUX_1024_1_IN_SEL = "1100000000" ELSE
				MUX_1024_1_IN_769 WHEN MUX_1024_1_IN_SEL = "1100000001" ELSE
				MUX_1024_1_IN_770 WHEN MUX_1024_1_IN_SEL = "1100000010" ELSE
				MUX_1024_1_IN_771 WHEN MUX_1024_1_IN_SEL = "1100000011" ELSE
				MUX_1024_1_IN_772 WHEN MUX_1024_1_IN_SEL = "1100000100" ELSE
				MUX_1024_1_IN_773 WHEN MUX_1024_1_IN_SEL = "1100000101" ELSE
				MUX_1024_1_IN_774 WHEN MUX_1024_1_IN_SEL = "1100000110" ELSE
				MUX_1024_1_IN_775 WHEN MUX_1024_1_IN_SEL = "1100000111" ELSE
				MUX_1024_1_IN_776 WHEN MUX_1024_1_IN_SEL = "1100001000" ELSE
				MUX_1024_1_IN_777 WHEN MUX_1024_1_IN_SEL = "1100001001" ELSE
				MUX_1024_1_IN_778 WHEN MUX_1024_1_IN_SEL = "1100001010" ELSE
				MUX_1024_1_IN_779 WHEN MUX_1024_1_IN_SEL = "1100001011" ELSE
				MUX_1024_1_IN_780 WHEN MUX_1024_1_IN_SEL = "1100001100" ELSE
				MUX_1024_1_IN_781 WHEN MUX_1024_1_IN_SEL = "1100001101" ELSE
				MUX_1024_1_IN_782 WHEN MUX_1024_1_IN_SEL = "1100001110" ELSE
				MUX_1024_1_IN_783 WHEN MUX_1024_1_IN_SEL = "1100001111" ELSE
				MUX_1024_1_IN_784 WHEN MUX_1024_1_IN_SEL = "1100010000" ELSE
				MUX_1024_1_IN_785 WHEN MUX_1024_1_IN_SEL = "1100010001" ELSE
				MUX_1024_1_IN_786 WHEN MUX_1024_1_IN_SEL = "1100010010" ELSE
				MUX_1024_1_IN_787 WHEN MUX_1024_1_IN_SEL = "1100010011" ELSE
				MUX_1024_1_IN_788 WHEN MUX_1024_1_IN_SEL = "1100010100" ELSE
				MUX_1024_1_IN_789 WHEN MUX_1024_1_IN_SEL = "1100010101" ELSE
				MUX_1024_1_IN_790 WHEN MUX_1024_1_IN_SEL = "1100010110" ELSE
				MUX_1024_1_IN_791 WHEN MUX_1024_1_IN_SEL = "1100010111" ELSE
				MUX_1024_1_IN_792 WHEN MUX_1024_1_IN_SEL = "1100011000" ELSE
				MUX_1024_1_IN_793 WHEN MUX_1024_1_IN_SEL = "1100011001" ELSE
				MUX_1024_1_IN_794 WHEN MUX_1024_1_IN_SEL = "1100011010" ELSE
				MUX_1024_1_IN_795 WHEN MUX_1024_1_IN_SEL = "1100011011" ELSE
				MUX_1024_1_IN_796 WHEN MUX_1024_1_IN_SEL = "1100011100" ELSE
				MUX_1024_1_IN_797 WHEN MUX_1024_1_IN_SEL = "1100011101" ELSE
				MUX_1024_1_IN_798 WHEN MUX_1024_1_IN_SEL = "1100011110" ELSE
				MUX_1024_1_IN_799 WHEN MUX_1024_1_IN_SEL = "1100011111" ELSE
				MUX_1024_1_IN_800 WHEN MUX_1024_1_IN_SEL = "1100100000" ELSE
				MUX_1024_1_IN_801 WHEN MUX_1024_1_IN_SEL = "1100100001" ELSE
				MUX_1024_1_IN_802 WHEN MUX_1024_1_IN_SEL = "1100100010" ELSE
				MUX_1024_1_IN_803 WHEN MUX_1024_1_IN_SEL = "1100100011" ELSE
				MUX_1024_1_IN_804 WHEN MUX_1024_1_IN_SEL = "1100100100" ELSE
				MUX_1024_1_IN_805 WHEN MUX_1024_1_IN_SEL = "1100100101" ELSE
				MUX_1024_1_IN_806 WHEN MUX_1024_1_IN_SEL = "1100100110" ELSE
				MUX_1024_1_IN_807 WHEN MUX_1024_1_IN_SEL = "1100100111" ELSE
				MUX_1024_1_IN_808 WHEN MUX_1024_1_IN_SEL = "1100101000" ELSE
				MUX_1024_1_IN_809 WHEN MUX_1024_1_IN_SEL = "1100101001" ELSE
				MUX_1024_1_IN_810 WHEN MUX_1024_1_IN_SEL = "1100101010" ELSE
				MUX_1024_1_IN_811 WHEN MUX_1024_1_IN_SEL = "1100101011" ELSE
				MUX_1024_1_IN_812 WHEN MUX_1024_1_IN_SEL = "1100101100" ELSE
				MUX_1024_1_IN_813 WHEN MUX_1024_1_IN_SEL = "1100101101" ELSE
				MUX_1024_1_IN_814 WHEN MUX_1024_1_IN_SEL = "1100101110" ELSE
				MUX_1024_1_IN_815 WHEN MUX_1024_1_IN_SEL = "1100101111" ELSE
				MUX_1024_1_IN_816 WHEN MUX_1024_1_IN_SEL = "1100110000" ELSE
				MUX_1024_1_IN_817 WHEN MUX_1024_1_IN_SEL = "1100110001" ELSE
				MUX_1024_1_IN_818 WHEN MUX_1024_1_IN_SEL = "1100110010" ELSE
				MUX_1024_1_IN_819 WHEN MUX_1024_1_IN_SEL = "1100110011" ELSE
				MUX_1024_1_IN_820 WHEN MUX_1024_1_IN_SEL = "1100110100" ELSE
				MUX_1024_1_IN_821 WHEN MUX_1024_1_IN_SEL = "1100110101" ELSE
				MUX_1024_1_IN_822 WHEN MUX_1024_1_IN_SEL = "1100110110" ELSE
				MUX_1024_1_IN_823 WHEN MUX_1024_1_IN_SEL = "1100110111" ELSE
				MUX_1024_1_IN_824 WHEN MUX_1024_1_IN_SEL = "1100111000" ELSE
				MUX_1024_1_IN_825 WHEN MUX_1024_1_IN_SEL = "1100111001" ELSE
				MUX_1024_1_IN_826 WHEN MUX_1024_1_IN_SEL = "1100111010" ELSE
				MUX_1024_1_IN_827 WHEN MUX_1024_1_IN_SEL = "1100111011" ELSE
				MUX_1024_1_IN_828 WHEN MUX_1024_1_IN_SEL = "1100111100" ELSE
				MUX_1024_1_IN_829 WHEN MUX_1024_1_IN_SEL = "1100111101" ELSE
				MUX_1024_1_IN_830 WHEN MUX_1024_1_IN_SEL = "1100111110" ELSE
				MUX_1024_1_IN_831 WHEN MUX_1024_1_IN_SEL = "1100111111" ELSE
				MUX_1024_1_IN_832 WHEN MUX_1024_1_IN_SEL = "1101000000" ELSE
				MUX_1024_1_IN_833 WHEN MUX_1024_1_IN_SEL = "1101000001" ELSE
				MUX_1024_1_IN_834 WHEN MUX_1024_1_IN_SEL = "1101000010" ELSE
				MUX_1024_1_IN_835 WHEN MUX_1024_1_IN_SEL = "1101000011" ELSE
				MUX_1024_1_IN_836 WHEN MUX_1024_1_IN_SEL = "1101000100" ELSE
				MUX_1024_1_IN_837 WHEN MUX_1024_1_IN_SEL = "1101000101" ELSE
				MUX_1024_1_IN_838 WHEN MUX_1024_1_IN_SEL = "1101000110" ELSE
				MUX_1024_1_IN_839 WHEN MUX_1024_1_IN_SEL = "1101000111" ELSE
				MUX_1024_1_IN_840 WHEN MUX_1024_1_IN_SEL = "1101001000" ELSE
				MUX_1024_1_IN_841 WHEN MUX_1024_1_IN_SEL = "1101001001" ELSE
				MUX_1024_1_IN_842 WHEN MUX_1024_1_IN_SEL = "1101001010" ELSE
				MUX_1024_1_IN_843 WHEN MUX_1024_1_IN_SEL = "1101001011" ELSE
				MUX_1024_1_IN_844 WHEN MUX_1024_1_IN_SEL = "1101001100" ELSE
				MUX_1024_1_IN_845 WHEN MUX_1024_1_IN_SEL = "1101001101" ELSE
				MUX_1024_1_IN_846 WHEN MUX_1024_1_IN_SEL = "1101001110" ELSE
				MUX_1024_1_IN_847 WHEN MUX_1024_1_IN_SEL = "1101001111" ELSE
				MUX_1024_1_IN_848 WHEN MUX_1024_1_IN_SEL = "1101010000" ELSE
				MUX_1024_1_IN_849 WHEN MUX_1024_1_IN_SEL = "1101010001" ELSE
				MUX_1024_1_IN_850 WHEN MUX_1024_1_IN_SEL = "1101010010" ELSE
				MUX_1024_1_IN_851 WHEN MUX_1024_1_IN_SEL = "1101010011" ELSE
				MUX_1024_1_IN_852 WHEN MUX_1024_1_IN_SEL = "1101010100" ELSE
				MUX_1024_1_IN_853 WHEN MUX_1024_1_IN_SEL = "1101010101" ELSE
				MUX_1024_1_IN_854 WHEN MUX_1024_1_IN_SEL = "1101010110" ELSE
				MUX_1024_1_IN_855 WHEN MUX_1024_1_IN_SEL = "1101010111" ELSE
				MUX_1024_1_IN_856 WHEN MUX_1024_1_IN_SEL = "1101011000" ELSE
				MUX_1024_1_IN_857 WHEN MUX_1024_1_IN_SEL = "1101011001" ELSE
				MUX_1024_1_IN_858 WHEN MUX_1024_1_IN_SEL = "1101011010" ELSE
				MUX_1024_1_IN_859 WHEN MUX_1024_1_IN_SEL = "1101011011" ELSE
				MUX_1024_1_IN_860 WHEN MUX_1024_1_IN_SEL = "1101011100" ELSE
				MUX_1024_1_IN_861 WHEN MUX_1024_1_IN_SEL = "1101011101" ELSE
				MUX_1024_1_IN_862 WHEN MUX_1024_1_IN_SEL = "1101011110" ELSE
				MUX_1024_1_IN_863 WHEN MUX_1024_1_IN_SEL = "1101011111" ELSE
				MUX_1024_1_IN_864 WHEN MUX_1024_1_IN_SEL = "1101100000" ELSE
				MUX_1024_1_IN_865 WHEN MUX_1024_1_IN_SEL = "1101100001" ELSE
				MUX_1024_1_IN_866 WHEN MUX_1024_1_IN_SEL = "1101100010" ELSE
				MUX_1024_1_IN_867 WHEN MUX_1024_1_IN_SEL = "1101100011" ELSE
				MUX_1024_1_IN_868 WHEN MUX_1024_1_IN_SEL = "1101100100" ELSE
				MUX_1024_1_IN_869 WHEN MUX_1024_1_IN_SEL = "1101100101" ELSE
				MUX_1024_1_IN_870 WHEN MUX_1024_1_IN_SEL = "1101100110" ELSE
				MUX_1024_1_IN_871 WHEN MUX_1024_1_IN_SEL = "1101100111" ELSE
				MUX_1024_1_IN_872 WHEN MUX_1024_1_IN_SEL = "1101101000" ELSE
				MUX_1024_1_IN_873 WHEN MUX_1024_1_IN_SEL = "1101101001" ELSE
				MUX_1024_1_IN_874 WHEN MUX_1024_1_IN_SEL = "1101101010" ELSE
				MUX_1024_1_IN_875 WHEN MUX_1024_1_IN_SEL = "1101101011" ELSE
				MUX_1024_1_IN_876 WHEN MUX_1024_1_IN_SEL = "1101101100" ELSE
				MUX_1024_1_IN_877 WHEN MUX_1024_1_IN_SEL = "1101101101" ELSE
				MUX_1024_1_IN_878 WHEN MUX_1024_1_IN_SEL = "1101101110" ELSE
				MUX_1024_1_IN_879 WHEN MUX_1024_1_IN_SEL = "1101101111" ELSE
				MUX_1024_1_IN_880 WHEN MUX_1024_1_IN_SEL = "1101110000" ELSE
				MUX_1024_1_IN_881 WHEN MUX_1024_1_IN_SEL = "1101110001" ELSE
				MUX_1024_1_IN_882 WHEN MUX_1024_1_IN_SEL = "1101110010" ELSE
				MUX_1024_1_IN_883 WHEN MUX_1024_1_IN_SEL = "1101110011" ELSE
				MUX_1024_1_IN_884 WHEN MUX_1024_1_IN_SEL = "1101110100" ELSE
				MUX_1024_1_IN_885 WHEN MUX_1024_1_IN_SEL = "1101110101" ELSE
				MUX_1024_1_IN_886 WHEN MUX_1024_1_IN_SEL = "1101110110" ELSE
				MUX_1024_1_IN_887 WHEN MUX_1024_1_IN_SEL = "1101110111" ELSE
				MUX_1024_1_IN_888 WHEN MUX_1024_1_IN_SEL = "1101111000" ELSE
				MUX_1024_1_IN_889 WHEN MUX_1024_1_IN_SEL = "1101111001" ELSE
				MUX_1024_1_IN_890 WHEN MUX_1024_1_IN_SEL = "1101111010" ELSE
				MUX_1024_1_IN_891 WHEN MUX_1024_1_IN_SEL = "1101111011" ELSE
				MUX_1024_1_IN_892 WHEN MUX_1024_1_IN_SEL = "1101111100" ELSE
				MUX_1024_1_IN_893 WHEN MUX_1024_1_IN_SEL = "1101111101" ELSE
				MUX_1024_1_IN_894 WHEN MUX_1024_1_IN_SEL = "1101111110" ELSE
				MUX_1024_1_IN_895 WHEN MUX_1024_1_IN_SEL = "1101111111" ELSE
				MUX_1024_1_IN_896 WHEN MUX_1024_1_IN_SEL = "1110000000" ELSE
				MUX_1024_1_IN_897 WHEN MUX_1024_1_IN_SEL = "1110000001" ELSE
				MUX_1024_1_IN_898 WHEN MUX_1024_1_IN_SEL = "1110000010" ELSE
				MUX_1024_1_IN_899 WHEN MUX_1024_1_IN_SEL = "1110000011" ELSE
				MUX_1024_1_IN_900 WHEN MUX_1024_1_IN_SEL = "1110000100" ELSE
				MUX_1024_1_IN_901 WHEN MUX_1024_1_IN_SEL = "1110000101" ELSE
				MUX_1024_1_IN_902 WHEN MUX_1024_1_IN_SEL = "1110000110" ELSE
				MUX_1024_1_IN_903 WHEN MUX_1024_1_IN_SEL = "1110000111" ELSE
				MUX_1024_1_IN_904 WHEN MUX_1024_1_IN_SEL = "1110001000" ELSE
				MUX_1024_1_IN_905 WHEN MUX_1024_1_IN_SEL = "1110001001" ELSE
				MUX_1024_1_IN_906 WHEN MUX_1024_1_IN_SEL = "1110001010" ELSE
				MUX_1024_1_IN_907 WHEN MUX_1024_1_IN_SEL = "1110001011" ELSE
				MUX_1024_1_IN_908 WHEN MUX_1024_1_IN_SEL = "1110001100" ELSE
				MUX_1024_1_IN_909 WHEN MUX_1024_1_IN_SEL = "1110001101" ELSE
				MUX_1024_1_IN_910 WHEN MUX_1024_1_IN_SEL = "1110001110" ELSE
				MUX_1024_1_IN_911 WHEN MUX_1024_1_IN_SEL = "1110001111" ELSE
				MUX_1024_1_IN_912 WHEN MUX_1024_1_IN_SEL = "1110010000" ELSE
				MUX_1024_1_IN_913 WHEN MUX_1024_1_IN_SEL = "1110010001" ELSE
				MUX_1024_1_IN_914 WHEN MUX_1024_1_IN_SEL = "1110010010" ELSE
				MUX_1024_1_IN_915 WHEN MUX_1024_1_IN_SEL = "1110010011" ELSE
				MUX_1024_1_IN_916 WHEN MUX_1024_1_IN_SEL = "1110010100" ELSE
				MUX_1024_1_IN_917 WHEN MUX_1024_1_IN_SEL = "1110010101" ELSE
				MUX_1024_1_IN_918 WHEN MUX_1024_1_IN_SEL = "1110010110" ELSE
				MUX_1024_1_IN_919 WHEN MUX_1024_1_IN_SEL = "1110010111" ELSE
				MUX_1024_1_IN_920 WHEN MUX_1024_1_IN_SEL = "1110011000" ELSE
				MUX_1024_1_IN_921 WHEN MUX_1024_1_IN_SEL = "1110011001" ELSE
				MUX_1024_1_IN_922 WHEN MUX_1024_1_IN_SEL = "1110011010" ELSE
				MUX_1024_1_IN_923 WHEN MUX_1024_1_IN_SEL = "1110011011" ELSE
				MUX_1024_1_IN_924 WHEN MUX_1024_1_IN_SEL = "1110011100" ELSE
				MUX_1024_1_IN_925 WHEN MUX_1024_1_IN_SEL = "1110011101" ELSE
				MUX_1024_1_IN_926 WHEN MUX_1024_1_IN_SEL = "1110011110" ELSE
				MUX_1024_1_IN_927 WHEN MUX_1024_1_IN_SEL = "1110011111" ELSE
				MUX_1024_1_IN_928 WHEN MUX_1024_1_IN_SEL = "1110100000" ELSE
				MUX_1024_1_IN_929 WHEN MUX_1024_1_IN_SEL = "1110100001" ELSE
				MUX_1024_1_IN_930 WHEN MUX_1024_1_IN_SEL = "1110100010" ELSE
				MUX_1024_1_IN_931 WHEN MUX_1024_1_IN_SEL = "1110100011" ELSE
				MUX_1024_1_IN_932 WHEN MUX_1024_1_IN_SEL = "1110100100" ELSE
				MUX_1024_1_IN_933 WHEN MUX_1024_1_IN_SEL = "1110100101" ELSE
				MUX_1024_1_IN_934 WHEN MUX_1024_1_IN_SEL = "1110100110" ELSE
				MUX_1024_1_IN_935 WHEN MUX_1024_1_IN_SEL = "1110100111" ELSE
				MUX_1024_1_IN_936 WHEN MUX_1024_1_IN_SEL = "1110101000" ELSE
				MUX_1024_1_IN_937 WHEN MUX_1024_1_IN_SEL = "1110101001" ELSE
				MUX_1024_1_IN_938 WHEN MUX_1024_1_IN_SEL = "1110101010" ELSE
				MUX_1024_1_IN_939 WHEN MUX_1024_1_IN_SEL = "1110101011" ELSE
				MUX_1024_1_IN_940 WHEN MUX_1024_1_IN_SEL = "1110101100" ELSE
				MUX_1024_1_IN_941 WHEN MUX_1024_1_IN_SEL = "1110101101" ELSE
				MUX_1024_1_IN_942 WHEN MUX_1024_1_IN_SEL = "1110101110" ELSE
				MUX_1024_1_IN_943 WHEN MUX_1024_1_IN_SEL = "1110101111" ELSE
				MUX_1024_1_IN_944 WHEN MUX_1024_1_IN_SEL = "1110110000" ELSE
				MUX_1024_1_IN_945 WHEN MUX_1024_1_IN_SEL = "1110110001" ELSE
				MUX_1024_1_IN_946 WHEN MUX_1024_1_IN_SEL = "1110110010" ELSE
				MUX_1024_1_IN_947 WHEN MUX_1024_1_IN_SEL = "1110110011" ELSE
				MUX_1024_1_IN_948 WHEN MUX_1024_1_IN_SEL = "1110110100" ELSE
				MUX_1024_1_IN_949 WHEN MUX_1024_1_IN_SEL = "1110110101" ELSE
				MUX_1024_1_IN_950 WHEN MUX_1024_1_IN_SEL = "1110110110" ELSE
				MUX_1024_1_IN_951 WHEN MUX_1024_1_IN_SEL = "1110110111" ELSE
				MUX_1024_1_IN_952 WHEN MUX_1024_1_IN_SEL = "1110111000" ELSE
				MUX_1024_1_IN_953 WHEN MUX_1024_1_IN_SEL = "1110111001" ELSE
				MUX_1024_1_IN_954 WHEN MUX_1024_1_IN_SEL = "1110111010" ELSE
				MUX_1024_1_IN_955 WHEN MUX_1024_1_IN_SEL = "1110111011" ELSE
				MUX_1024_1_IN_956 WHEN MUX_1024_1_IN_SEL = "1110111100" ELSE
				MUX_1024_1_IN_957 WHEN MUX_1024_1_IN_SEL = "1110111101" ELSE
				MUX_1024_1_IN_958 WHEN MUX_1024_1_IN_SEL = "1110111110" ELSE
				MUX_1024_1_IN_959 WHEN MUX_1024_1_IN_SEL = "1110111111" ELSE
				MUX_1024_1_IN_960 WHEN MUX_1024_1_IN_SEL = "1111000000" ELSE
				MUX_1024_1_IN_961 WHEN MUX_1024_1_IN_SEL = "1111000001" ELSE
				MUX_1024_1_IN_962 WHEN MUX_1024_1_IN_SEL = "1111000010" ELSE
				MUX_1024_1_IN_963 WHEN MUX_1024_1_IN_SEL = "1111000011" ELSE
				MUX_1024_1_IN_964 WHEN MUX_1024_1_IN_SEL = "1111000100" ELSE
				MUX_1024_1_IN_965 WHEN MUX_1024_1_IN_SEL = "1111000101" ELSE
				MUX_1024_1_IN_966 WHEN MUX_1024_1_IN_SEL = "1111000110" ELSE
				MUX_1024_1_IN_967 WHEN MUX_1024_1_IN_SEL = "1111000111" ELSE
				MUX_1024_1_IN_968 WHEN MUX_1024_1_IN_SEL = "1111001000" ELSE
				MUX_1024_1_IN_969 WHEN MUX_1024_1_IN_SEL = "1111001001" ELSE
				MUX_1024_1_IN_970 WHEN MUX_1024_1_IN_SEL = "1111001010" ELSE
				MUX_1024_1_IN_971 WHEN MUX_1024_1_IN_SEL = "1111001011" ELSE
				MUX_1024_1_IN_972 WHEN MUX_1024_1_IN_SEL = "1111001100" ELSE
				MUX_1024_1_IN_973 WHEN MUX_1024_1_IN_SEL = "1111001101" ELSE
				MUX_1024_1_IN_974 WHEN MUX_1024_1_IN_SEL = "1111001110" ELSE
				MUX_1024_1_IN_975 WHEN MUX_1024_1_IN_SEL = "1111001111" ELSE
				MUX_1024_1_IN_976 WHEN MUX_1024_1_IN_SEL = "1111010000" ELSE
				MUX_1024_1_IN_977 WHEN MUX_1024_1_IN_SEL = "1111010001" ELSE
				MUX_1024_1_IN_978 WHEN MUX_1024_1_IN_SEL = "1111010010" ELSE
				MUX_1024_1_IN_979 WHEN MUX_1024_1_IN_SEL = "1111010011" ELSE
				MUX_1024_1_IN_980 WHEN MUX_1024_1_IN_SEL = "1111010100" ELSE
				MUX_1024_1_IN_981 WHEN MUX_1024_1_IN_SEL = "1111010101" ELSE
				MUX_1024_1_IN_982 WHEN MUX_1024_1_IN_SEL = "1111010110" ELSE
				MUX_1024_1_IN_983 WHEN MUX_1024_1_IN_SEL = "1111010111" ELSE
				MUX_1024_1_IN_984 WHEN MUX_1024_1_IN_SEL = "1111011000" ELSE
				MUX_1024_1_IN_985 WHEN MUX_1024_1_IN_SEL = "1111011001" ELSE
				MUX_1024_1_IN_986 WHEN MUX_1024_1_IN_SEL = "1111011010" ELSE
				MUX_1024_1_IN_987 WHEN MUX_1024_1_IN_SEL = "1111011011" ELSE
				MUX_1024_1_IN_988 WHEN MUX_1024_1_IN_SEL = "1111011100" ELSE
				MUX_1024_1_IN_989 WHEN MUX_1024_1_IN_SEL = "1111011101" ELSE
				MUX_1024_1_IN_990 WHEN MUX_1024_1_IN_SEL = "1111011110" ELSE
				MUX_1024_1_IN_991 WHEN MUX_1024_1_IN_SEL = "1111011111" ELSE
				MUX_1024_1_IN_992 WHEN MUX_1024_1_IN_SEL = "1111100000" ELSE
				MUX_1024_1_IN_993 WHEN MUX_1024_1_IN_SEL = "1111100001" ELSE
				MUX_1024_1_IN_994 WHEN MUX_1024_1_IN_SEL = "1111100010" ELSE
				MUX_1024_1_IN_995 WHEN MUX_1024_1_IN_SEL = "1111100011" ELSE
				MUX_1024_1_IN_996 WHEN MUX_1024_1_IN_SEL = "1111100100" ELSE
				MUX_1024_1_IN_997 WHEN MUX_1024_1_IN_SEL = "1111100101" ELSE
				MUX_1024_1_IN_998 WHEN MUX_1024_1_IN_SEL = "1111100110" ELSE
				MUX_1024_1_IN_999 WHEN MUX_1024_1_IN_SEL = "1111100111" ELSE
				MUX_1024_1_IN_1000 WHEN MUX_1024_1_IN_SEL = "1111101000" ELSE
				MUX_1024_1_IN_1001 WHEN MUX_1024_1_IN_SEL = "1111101001" ELSE
				MUX_1024_1_IN_1002 WHEN MUX_1024_1_IN_SEL = "1111101010" ELSE
				MUX_1024_1_IN_1003 WHEN MUX_1024_1_IN_SEL = "1111101011" ELSE
				MUX_1024_1_IN_1004 WHEN MUX_1024_1_IN_SEL = "1111101100" ELSE
				MUX_1024_1_IN_1005 WHEN MUX_1024_1_IN_SEL = "1111101101" ELSE
				MUX_1024_1_IN_1006 WHEN MUX_1024_1_IN_SEL = "1111101110" ELSE
				MUX_1024_1_IN_1007 WHEN MUX_1024_1_IN_SEL = "1111101111" ELSE
				MUX_1024_1_IN_1008 WHEN MUX_1024_1_IN_SEL = "1111110000" ELSE
				MUX_1024_1_IN_1009 WHEN MUX_1024_1_IN_SEL = "1111110001" ELSE
				MUX_1024_1_IN_1010 WHEN MUX_1024_1_IN_SEL = "1111110010" ELSE
				MUX_1024_1_IN_1011 WHEN MUX_1024_1_IN_SEL = "1111110011" ELSE
				MUX_1024_1_IN_1012 WHEN MUX_1024_1_IN_SEL = "1111110100" ELSE
				MUX_1024_1_IN_1013 WHEN MUX_1024_1_IN_SEL = "1111110101" ELSE
				MUX_1024_1_IN_1014 WHEN MUX_1024_1_IN_SEL = "1111110110" ELSE
				MUX_1024_1_IN_1015 WHEN MUX_1024_1_IN_SEL = "1111110111" ELSE
				MUX_1024_1_IN_1016 WHEN MUX_1024_1_IN_SEL = "1111111000" ELSE
				MUX_1024_1_IN_1017 WHEN MUX_1024_1_IN_SEL = "1111111001" ELSE
				MUX_1024_1_IN_1018 WHEN MUX_1024_1_IN_SEL = "1111111010" ELSE
				MUX_1024_1_IN_1019 WHEN MUX_1024_1_IN_SEL = "1111111011" ELSE
				MUX_1024_1_IN_1020 WHEN MUX_1024_1_IN_SEL = "1111111100" ELSE
				MUX_1024_1_IN_1021 WHEN MUX_1024_1_IN_SEL = "1111111101" ELSE
				MUX_1024_1_IN_1022 WHEN MUX_1024_1_IN_SEL = "1111111110" ELSE
				MUX_1024_1_IN_1023 WHEN MUX_1024_1_IN_SEL = "1111111111" ELSE
				(OTHERS => '0');


END behavioral;