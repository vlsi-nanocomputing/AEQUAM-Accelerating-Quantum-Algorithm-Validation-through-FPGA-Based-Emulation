LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EMULATOR_N_6_W_2_S_0_Q_2 IS
GENERIC( K : INTEGER := 20 );
PORT (
	EMULATOR_N_6_W_2_S_0_Q_2_IN_FROM_MCU : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
	EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK : IN STD_LOGIC;
	EMULATOR_N_6_W_2_S_0_Q_2_IN_RSTN : IN STD_LOGIC;
	EMULATOR_N_6_W_2_S_0_Q_2_OUT_TO_MCU : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
	EMULATOR_N_6_W_2_S_0_Q_2_IN_OUT_BUS : INOUT STD_LOGIC_VECTOR (K-1 DOWNTO 0)
);
END ENTITY;
ARCHITECTURE generated OF EMULATOR_N_6_W_2_S_0_Q_2 IS
COMPONENT QPE_control IS
PORT (
		QPE_CONTROL_IN_FROM_MCU : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		QPE_CONTROL_IN_ACK : IN STD_LOGIC;
		QPE_CONTROL_IN_COMPLETED : IN STD_LOGIC;
      QPE_CONTROL_IN_GATE_COMP : IN STD_LOGIC;
		QPE_CONTROL_IN_CLK : IN STD_LOGIC;
        QPE_CONTROL_IN_RSTN : IN STD_LOGIC;
		QPE_CONTROL_OUT_TO_MCU : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		QPE_CONTROL_OUT_CLR_ALL : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAVE_QUBIT_NUMB : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAMPLE_INSTR : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAMPLE_SIN_COS : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAVE_SIN_COS : OUT STD_LOGIC;
		QPE_CONTROL_OUT_EN_RES_CNT : OUT STD_LOGIC;
       QPE_CONTROL_OUT_EN_OUT_BUF : OUT STD_LOGIC;
       QPE_CONTROL_OUT_MCU_ACK_TOGGLE : OUT STD_LOGIC;
QPE_CONTROL_OUT_EN_QEP_DONE : OUT STD_LOGIC
	);
END COMPONENT;
COMPONENT counter IS
GENERIC (N : NATURAL := 32);
PORT (
COUNTER_IN_EN : IN STD_LOGIC;
COUNTER_IN_CLR : IN STD_LOGIC;
COUNTER_IN_CLK : IN STD_LOGIC;
COUNTER_OUT_DATA : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END COMPONENT;COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_2_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_2_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		MUX_2_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_4_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_4_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_4_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_4_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_4_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_4_1_IN_SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		MUX_4_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT state_decoder_N_6 IS
 PORT (
 STATE_DECODER_N_6_IN_QTGT : IN STD_LOGIC_VECTOR( 2 DOWNTO 0);
 STATE_DECODER_N_6_IN_QCTRL : IN STD_LOGIC_VECTOR( 2 DOWNTO 0);
 STATE_DECODER_N_6_IN_OPCODE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
 STATE_DECODER_N_6_IN_SAVE_QBIT_NUMBER : IN STD_LOGIC;
 STATE_DECODER_N_6_IN_CLEAR : IN STD_LOGIC;
 STATE_DECODER_N_6_IN_CLK : IN STD_LOGIC;
 STATE_DECODER_N_6_OUT_MASK_FIRST : OUT STD_LOGIC;  
STATE_DECODER_N_6_OUT_CTRL_MASK : OUT STD_LOGIC_VECTOR ( 63 DOWNTO 0)
 );
 END COMPONENT;
COMPONENT QEP_N_6_W_2_S_0 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		QEP_N_6_W_2_S_0_IN_START : IN STD_LOGIC;
		QEP_N_6_W_2_S_0_IN_QTGT : IN STD_LOGIC_VECTOR (2 DOWNTO 0); 
		QEP_N_6_W_2_S_0_IN_CTRL_MASK : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		QEP_N_6_W_2_S_0_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		QEP_N_6_W_2_S_0_IN_SIN : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_6_W_2_S_0_IN_COS : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_6_W_2_S_0_IN_WIN_SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		QEP_N_6_W_2_S_0_IN_OUT_STATE_SEL : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		QEP_N_6_W_2_S_0_IN_REAL_IMAG_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		QEP_N_6_W_2_S_0_IN_CLK : IN STD_LOGIC;
		QEP_N_6_W_2_S_0_IN_CLEAR : IN STD_LOGIC;
		QEP_N_6_W_2_S_0_IN_MASK_FIRST_COEFF : IN STD_LOGIC;
		QEP_N_6_W_2_S_0_IN_ENABLE_STATE_UPDATE : IN STD_LOGIC;
		QEP_N_6_W_2_S_0_OUT_DONE : OUT STD_LOGIC;
		QEP_N_6_W_2_S_0_OUT_DATA : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT
;SIGNAL FROM_QPE_CTRL_EN_QEP_DONE, GATE_COMPLETE, FETCH_INSTRUCTION, TO_QPE_CTRL_ACK, TO_QPE_CTRL_COMPLETE, FROM_QPE_CTRL_SAMPLE_SIN_COS, FROM_QPE_CTRL_SAVE_SIN_COS, FROM_QPE_CTRL_CLEAR, FROM_QPE_CTRL_SAMPLE_INSTR, FROM_QPE_CTRL_SAVE_QBIT_NUMB, FROM_QPE_CTRL_EN_RES_CNT : STD_LOGIC;
SIGNAL FROM_TRIG_ADD_SIN_COS_ADD : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL FROM_DEC_MASK_FIRST : STD_LOGIC;
SIGNAL FROM_DEC_QIMM : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL FROM_TRIG_UNIT_SIN, FROM_TRIG_UNIT_COS, FROM_FETCH_SIN_COS : STD_LOGIC_VECTOR (K-1 DOWNTO 0);SIGNAL ROW_SEL_SIN_COS, ENABLE_SIN_DEC, ENABLE_COS_DEC : STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL FROM_SIN_REG_0,FROM_SIN_REG_1,FROM_SIN_REG_2,FROM_SIN_REG_3: STD_LOGIC_VECTOR(K-1 DOWNTO 0);
SIGNAL FROM_COS_REG_0,FROM_COS_REG_1,FROM_COS_REG_2,FROM_COS_REG_3: STD_LOGIC_VECTOR(K-1 DOWNTO 0);
SIGNAL ENABLE_SIN_REG, ENABLE_COS_REG : STD_LOGIC;
SIGNAL FROM_FETCH_INSTR : STD_LOGIC_VECTOR(11 DOWNTO 0);SIGNAL CTRL_MASK : STD_LOGIC_VECTOR ( 63 DOWNTO 0);
SIGNAL OPCODE : STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL QTGT, QCTRL : STD_LOGIC_VECTOR (2 DOWNTO 0);
SIGNAL FROM_QEP_DONE, QEP_DONE_ENABLED, TO_QEP_START, TO_QEP_START_PIPE :STD_LOGIC;
SIGNAL FROM_WIN_CNT_TC : STD_LOGIC;
SIGNAL WINDOW_SELECTOR : STD_LOGIC_VECTOR( 1 DOWNTO 0);
SIGNAL RESULT_SELECTOR : STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL BUFFER_IN, BUFFER_OUT, RESULT : STD_LOGIC_VECTOR(K-1 DOWNTO 0);
SIGNAL OUT_BUF_EN, MCU_ACK_TOGGLE : STD_LOGIC;
BEGIN
QPE_CTRL: QPE_control PORT MAP(
		QPE_CONTROL_IN_FROM_MCU => EMULATOR_N_6_W_2_S_0_Q_2_IN_FROM_MCU ,
		QPE_CONTROL_IN_ACK => TO_QPE_CTRL_ACK ,
		QPE_CONTROL_IN_COMPLETED => TO_QPE_CTRL_COMPLETE , 
       QPE_CONTROL_IN_GATE_COMP => GATE_COMPLETE,
		QPE_CONTROL_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
     QPE_CONTROL_IN_RSTN => EMULATOR_N_6_W_2_S_0_Q_2_IN_RSTN,
		QPE_CONTROL_OUT_TO_MCU => EMULATOR_N_6_W_2_S_0_Q_2_OUT_TO_MCU ,
		QPE_CONTROL_OUT_CLR_ALL => FROM_QPE_CTRL_CLEAR ,
		QPE_CONTROL_OUT_SAVE_QUBIT_NUMB => FROM_QPE_CTRL_SAVE_QBIT_NUMB ,
		QPE_CONTROL_OUT_SAMPLE_INSTR => FROM_QPE_CTRL_SAMPLE_INSTR ,
		QPE_CONTROL_OUT_SAMPLE_SIN_COS => FROM_QPE_CTRL_SAMPLE_SIN_COS ,
		QPE_CONTROL_OUT_SAVE_SIN_COS => FROM_QPE_CTRL_SAVE_SIN_COS ,
		QPE_CONTROL_OUT_EN_RES_CNT => FROM_QPE_CTRL_EN_RES_CNT,
     QPE_CONTROL_OUT_EN_OUT_BUF => OUT_BUF_EN,
     QPE_CONTROL_OUT_MCU_ACK_TOGGLE => MCU_ACK_TOGGLE,
QPE_CONTROL_OUT_EN_QEP_DONE =>	FROM_QPE_CTRL_EN_QEP_DONE);
CNT_TRIG_ADD : counter GENERIC MAP (3)
PORT MAP (
COUNTER_IN_EN => FROM_QPE_CTRL_SAVE_SIN_COS ,
COUNTER_IN_CLR => FROM_QPE_CTRL_CLEAR,
COUNTER_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK,
COUNTER_OUT_DATA => FROM_TRIG_ADD_SIN_COS_ADD);
ENABLE_SIN_REG <= FROM_QPE_CTRL_SAVE_SIN_COS AND ( NOT FROM_TRIG_ADD_SIN_COS_ADD(0) );
ENABLE_COS_REG <= FROM_QPE_CTRL_SAVE_SIN_COS AND FROM_TRIG_ADD_SIN_COS_ADD(0);
ROW_SEL_SIN_COS <= 
"0001" WHEN FROM_TRIG_ADD_SIN_COS_ADD( 2 DOWNTO 1) = "00" ELSE
"0010" WHEN FROM_TRIG_ADD_SIN_COS_ADD( 2 DOWNTO 1) = "01" ELSE
"0100" WHEN FROM_TRIG_ADD_SIN_COS_ADD( 2 DOWNTO 1) = "10" ELSE
"1000" WHEN FROM_TRIG_ADD_SIN_COS_ADD( 2 DOWNTO 1) = "11" ELSE
(OTHERS => '0');
ENABLE_SIN_DEC(0) <= ENABLE_SIN_REG AND ROW_SEL_SIN_COS(0);
ENABLE_COS_DEC(0) <= ENABLE_COS_REG AND ROW_SEL_SIN_COS(0);
ENABLE_SIN_DEC(1) <= ENABLE_SIN_REG AND ROW_SEL_SIN_COS(1);
ENABLE_COS_DEC(1) <= ENABLE_COS_REG AND ROW_SEL_SIN_COS(1);
ENABLE_SIN_DEC(2) <= ENABLE_SIN_REG AND ROW_SEL_SIN_COS(2);
ENABLE_COS_DEC(2) <= ENABLE_COS_REG AND ROW_SEL_SIN_COS(2);
ENABLE_SIN_DEC(3) <= ENABLE_SIN_REG AND ROW_SEL_SIN_COS(3);
ENABLE_COS_DEC(3) <= ENABLE_COS_REG AND ROW_SEL_SIN_COS(3);
SIN_REG_0 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_SIN_DEC(0) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_SIN_REG_0);
COS_REG_0 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_COS_DEC(0) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_COS_REG_0);
SIN_REG_1 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_SIN_DEC(1) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_SIN_REG_1);
COS_REG_1 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_COS_DEC(1) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_COS_REG_1);
SIN_REG_2 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_SIN_DEC(2) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_SIN_REG_2);
COS_REG_2 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_COS_DEC(2) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_COS_REG_2);
SIN_REG_3 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_SIN_DEC(3) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_SIN_REG_3);
COS_REG_3 : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => FROM_FETCH_SIN_COS ,
												REG_IN_ENABLE => ENABLE_COS_DEC(3) ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_COS_REG_3);
SIN_SELECTION : multiplexer_4_1 	GENERIC MAP (K)
									PORT MAP (
										MUX_4_1_IN_0 => FROM_SIN_REG_0 ,
										MUX_4_1_IN_1 => FROM_SIN_REG_1 ,
										MUX_4_1_IN_2 => FROM_SIN_REG_2 ,
										MUX_4_1_IN_3 => FROM_SIN_REG_3 ,
				                    			MUX_4_1_IN_SEL => FROM_DEC_QIMM ,
										MUX_4_1_OUT_RES => FROM_TRIG_UNIT_SIN
									);
COS_SELECTION : multiplexer_4_1 	GENERIC MAP (K)
									PORT MAP (
										MUX_4_1_IN_0 => FROM_COS_REG_0 ,
										MUX_4_1_IN_1 => FROM_COS_REG_1 ,
										MUX_4_1_IN_2 => FROM_COS_REG_2 ,
										MUX_4_1_IN_3 => FROM_COS_REG_3 ,
				                    			MUX_4_1_IN_SEL => FROM_DEC_QIMM ,
										MUX_4_1_OUT_RES => FROM_TRIG_UNIT_COS
									);
BUFFER_IN <= EMULATOR_N_6_W_2_S_0_Q_2_IN_OUT_BUS;
REG_FETCH_SIN_COS : n_bit_register
GENERIC MAP (K)
PORT MAP(
												REG_IN_DATA => BUFFER_IN ,
												REG_IN_ENABLE => FROM_QPE_CTRL_SAMPLE_SIN_COS ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_FETCH_SIN_COS);
FETCH_INSTRUCTION <= FROM_QPE_CTRL_SAMPLE_INSTR;
TO_QPE_CTRL_ACK <= FROM_QPE_CTRL_SAMPLE_SIN_COS OR FETCH_INSTRUCTION;
REG_FETCH_INSTR : n_bit_register
GENERIC MAP (12)
PORT MAP(
												REG_IN_DATA => BUFFER_IN(11 DOWNTO 0) ,
												REG_IN_ENABLE => FETCH_INSTRUCTION ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA => FROM_FETCH_INSTR);
DEC_STAGE : state_decoder_N_6 
 PORT MAP (
 STATE_DECODER_N_6_IN_QTGT => QTGT,
 STATE_DECODER_N_6_IN_QCTRL => FROM_FETCH_INSTR( 4 DOWNTO 2),
 STATE_DECODER_N_6_IN_OPCODE => FROM_FETCH_INSTR(11 DOWNTO 8),
 STATE_DECODER_N_6_IN_SAVE_QBIT_NUMBER => FROM_QPE_CTRL_SAVE_QBIT_NUMB,
 STATE_DECODER_N_6_IN_CLEAR => FROM_QPE_CTRL_CLEAR,
 STATE_DECODER_N_6_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK,
 STATE_DECODER_N_6_OUT_MASK_FIRST => FROM_DEC_MASK_FIRST, 
STATE_DECODER_N_6_OUT_CTRL_MASK => CTRL_MASK
 );
FROM_DEC_QIMM <= FROM_FETCH_INSTR (1 DOWNTO 0);
OPCODE <= FROM_FETCH_INSTR(11 DOWNTO 8);
QTGT <= FROM_FETCH_INSTR(7 DOWNTO 5);
QEP_DONE_ENABLED <= FROM_QPE_CTRL_EN_QEP_DONE AND FROM_QEP_DONE;
CNT_WIN_SEL : counter GENERIC MAP (2)
PORT MAP (
COUNTER_IN_EN => QEP_DONE_ENABLED ,
COUNTER_IN_CLR => FROM_QPE_CTRL_CLEAR,
COUNTER_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK,
COUNTER_OUT_DATA => WINDOW_SELECTOR);
FROM_WIN_CNT_TC <= '1' WHEN WINDOW_SELECTOR = "11" ELSE '0';
GATE_COMPLETE <= FROM_WIN_CNT_TC AND FROM_QEP_DONE AND QEP_DONE_ENABLED;
CNT_RES_SEL : counter GENERIC MAP (7)
PORT MAP (
COUNTER_IN_EN => FROM_QPE_CTRL_EN_RES_CNT ,
COUNTER_IN_CLR => FROM_QPE_CTRL_CLEAR,
COUNTER_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK,
COUNTER_OUT_DATA => RESULT_SELECTOR);
TO_QPE_CTRL_COMPLETE <= '1' WHEN RESULT_SELECTOR = "1111111" ELSE '0';
TO_QEP_START_PIPE <= FETCH_INSTRUCTION AND NOT FROM_QPE_CTRL_SAVE_QBIT_NUMB;
REG_START_PIPE : n_bit_register
GENERIC MAP (1)
PORT MAP(
												REG_IN_DATA(0) => TO_QEP_START_PIPE ,
												REG_IN_ENABLE => '1' ,
												REG_IN_CLEAR => FROM_QPE_CTRL_CLEAR ,
												REG_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK ,
												REG_OUT_DATA(0) => TO_QEP_START);
QEP_UNIT : QEP_N_6_W_2_S_0 
	GENERIC MAP (K)
	PORT MAP (
		QEP_N_6_W_2_S_0_IN_START => TO_QEP_START,
		QEP_N_6_W_2_S_0_IN_QTGT => QTGT, 
		QEP_N_6_W_2_S_0_IN_CTRL_MASK => CTRL_MASK,
		QEP_N_6_W_2_S_0_IN_OPCODE => OPCODE,
		QEP_N_6_W_2_S_0_IN_SIN => FROM_TRIG_UNIT_SIN,
		QEP_N_6_W_2_S_0_IN_COS => FROM_TRIG_UNIT_COS ,
		QEP_N_6_W_2_S_0_IN_WIN_SEL => WINDOW_SELECTOR ,
		QEP_N_6_W_2_S_0_IN_OUT_STATE_SEL => RESULT_SELECTOR(6 DOWNTO 1) ,
		QEP_N_6_W_2_S_0_IN_REAL_IMAG_SEL => RESULT_SELECTOR(0 DOWNTO 0),
		QEP_N_6_W_2_S_0_IN_CLK => EMULATOR_N_6_W_2_S_0_Q_2_IN_CLK,
		QEP_N_6_W_2_S_0_IN_CLEAR  => FROM_QPE_CTRL_CLEAR,
		QEP_N_6_W_2_S_0_IN_MASK_FIRST_COEFF => FROM_DEC_MASK_FIRST,
		QEP_N_6_W_2_S_0_IN_ENABLE_STATE_UPDATE => FROM_QPE_CTRL_EN_QEP_DONE,
		QEP_N_6_W_2_S_0_OUT_DONE => FROM_QEP_DONE,
		QEP_N_6_W_2_S_0_OUT_DATA => RESULT);
BUFFER_OUT <= RESULT WHEN OUT_BUF_EN = '1' ELSE (OTHERS => 'Z');
EMULATOR_N_6_W_2_S_0_Q_2_IN_OUT_BUS <= BUFFER_OUT;
END generated;
