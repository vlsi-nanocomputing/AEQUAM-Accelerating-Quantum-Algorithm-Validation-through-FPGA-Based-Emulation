library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY adder_subtractor IS 
	GENERIC ( K : INTEGER := 20);
	PORT(
		ADD_SUB_IN_A : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		ADD_SUB_IN_B : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		ADD_SUB_IN_SUB : IN STD_LOGIC;
		ADD_SUB_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE chosen OF adder_subtractor IS

	COMPONENT comb_adder IS
	GENERIC( K : INTEGER := 20);
	PORT(
		COMB_ADD_IN_A : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		COMB_ADD_IN_B : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		COMB_ADD_IN_CIN : IN STD_LOGIC;
		
		COMB_ADD_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
	END COMPONENT;

	SIGNAL XOR_IN_B : STD_LOGIC_VECTOR(K-1 DOWNTO 0);

	--CHOOSE ADDER ARCHITECTURE
	FOR ALL: comb_adder USE ENTITY WORK.comb_adder(behavioral);

BEGIN

	XOR_BITWISE: FOR INDEX_XOR IN 0 TO K-1 GENERATE
	BEGIN
		XOR_IN_B(INDEX_XOR) <= ADD_SUB_IN_B(INDEX_XOR) XOR ADD_SUB_IN_SUB;
	END GENERATE XOR_BITWISE;

	ADDER: comb_adder 	GENERIC MAP(K => K)
						PORT MAP (
							COMB_ADD_IN_A => ADD_SUB_IN_A,
							COMB_ADD_IN_B => XOR_IN_B,
							COMB_ADD_IN_CIN => ADD_SUB_IN_SUB,
							COMB_ADD_OUT_RES => ADD_SUB_OUT_RES
						);

END chosen;