LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY counter IS
GENERIC (N : NATURAL := 32);
PORT (
COUNTER_IN_EN : IN STD_LOGIC;
COUNTER_IN_CLR : IN STD_LOGIC;
COUNTER_IN_CLK : IN STD_LOGIC;
COUNTER_OUT_DATA : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END COUNTER;

ARCHITECTURE behavioral OF counter IS
BEGIN
		CNT: PROCESS(COUNTER_IN_CLK)
			VARIABLE CNT : UNSIGNED(N-1 DOWNTO 0) := (OTHERS => '0'); 
			BEGIN
				IF (COUNTER_IN_CLK'EVENT AND COUNTER_IN_CLK = '1') THEN
					IF (COUNTER_IN_CLR = '1') THEN
						CNT := (OTHERS => '0');
					ELSE
						IF (COUNTER_IN_EN = '1') THEN
							CNT := CNT + 1;
						END IF;
					END IF;
					COUNTER_OUT_DATA <= STD_LOGIC_VECTOR(CNT);
				END IF;
		END PROCESS;
END behavioral;
