LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY QPE_control IS 
	PORT (
		QPE_CONTROL_IN_FROM_MCU : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		
		QPE_CONTROL_IN_ACK : IN STD_LOGIC;
		QPE_CONTROL_IN_COMPLETED : IN STD_LOGIC;
		QPE_CONTROL_IN_GATE_COMP : IN STD_LOGIC;
		
		QPE_CONTROL_IN_CLK : IN STD_LOGIC;
		QPE_CONTROL_IN_RSTN : IN STD_LOGIC;
		
		QPE_CONTROL_OUT_TO_MCU : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		
		QPE_CONTROL_OUT_CLR_ALL : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAVE_QUBIT_NUMB : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAMPLE_INSTR : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAMPLE_SIN_COS : OUT STD_LOGIC;
		QPE_CONTROL_OUT_SAVE_SIN_COS : OUT STD_LOGIC;
		QPE_CONTROL_OUT_EN_RES_CNT : OUT STD_LOGIC;
		QPE_CONTROL_OUT_EN_OUT_BUF : OUT STD_LOGIC;
		QPE_CONTROL_OUT_MCU_ACK_TOGGLE : OUT STD_LOGIC;
		QPE_CONTROL_OUT_EN_QEP_DONE : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE state_machine OF QPE_control IS 

	COMPONENT n_bit_register IS
		generic (n_bit: INTEGER);
		port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
				REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
				REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
	END COMPONENT;

	TYPE STATE_TYPE IS (RESET, INIT_0, INIT_0_IDLE, INIT_0_END, INIT_I, INIT_I_IDLE, INIT_I_END, INIT_II, INIT_II_IDLE, INIT_II_END, INIT_III, INIT_III_IDLE, INIT_III_END, START_I, START_I_IDLE, START_I_END, START_I_EXE, START_II, START_II_END, START_II_IDLE, START_II_EXE, SEND, SEND_IDLE, SEND_END);
	SIGNAL CURRENT_STATE : STATE_TYPE;

	SIGNAL CLR,RES_EN, ACK_INIT, DEL_ACK_FROM_QEP, CLR_GATE_COMP, SAVED_GATE_COMP : STD_LOGIC;
	--SIGNAL TO_MCU_TOGGLE, FROM_MCU_TOGGLE : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL FROM_MCU_ACK, MCU_ACK_TOGGLE : STD_LOGIC_VECTOR(0 DOWNTO 0);

BEGIN

	--TO_MCU_TOGGLE(0) <= FROM_MCU_TOGGLE(0) XOR (QPE_CONTROL_IN_ACK OR ACK_INIT);
	--TO_MCU_TOGGLE(1) <= FROM_MCU_TOGGLE(1) XOR RES_EN;
	

	REG_GATE_COMP : n_bit_register 		GENERIC MAP (1)
											PORT MAP (
												REG_IN_DATA => "1",
												REG_IN_ENABLE => QPE_CONTROL_IN_GATE_COMP ,
												REG_IN_CLEAR => CLR_GATE_COMP ,
												REG_IN_CLK => QPE_CONTROL_IN_CLK ,
												REG_OUT_DATA(0) => SAVED_GATE_COMP
											);

	--QPE_CONTROL_OUT_TO_MCU <= FROM_MCU_TOGGLE;

	REG_HAND_MCU : n_bit_register 		GENERIC MAP (1)
											PORT MAP (
												REG_IN_DATA(0) => QPE_CONTROL_IN_ACK ,
												REG_IN_ENABLE => '1' ,
												REG_IN_CLEAR => CLR ,
												REG_IN_CLK => QPE_CONTROL_IN_CLK ,
												REG_OUT_DATA(0) => DEL_ACK_FROM_QEP
											);
	MCU_ACK_TOGGLE(0) <= (FROM_MCU_ACK(0) XOR QPE_CONTROL_IN_FROM_MCU(0)) AND (NOT CLR);


	REG_FROM_MCU: n_bit_register		GENERIC MAP	(1)
											PORT MAP(
												REG_IN_DATA => QPE_CONTROL_IN_FROM_MCU(0 DOWNTO 0) ,
												REG_IN_ENABLE => '1' ,
												REG_IN_CLEAR => CLR ,
												REG_IN_CLK => QPE_CONTROL_IN_CLK ,
												REG_OUT_DATA => FROM_MCU_ACK
											);

	REG_DELAY_MCU_ACK: n_bit_register		GENERIC MAP	(1)
											PORT MAP(
												REG_IN_DATA => "1" ,
												REG_IN_ENABLE => MCU_ACK_TOGGLE(0) ,
												REG_IN_CLEAR => QPE_CONTROL_IN_ACK ,
												REG_IN_CLK => QPE_CONTROL_IN_CLK ,
												REG_OUT_DATA(0) => QPE_CONTROL_OUT_MCU_ACK_TOGGLE
											);
	
	--To MCU
	--TO_MCU : PROCESS (QPE_CONTROL_IN_CLK)
	--BEGIN
	
	--	IF RISING_EDGE(QPE_CONTROL_IN_CLK) THEN
		
	--		IF CLR <= '1' THEN
	--			PREV_ACK <= '0';
	--			PREV_READ <= '0';
	--		ELSE 
	--			PREV_ACK <= PREV_ACK XOR QPE_CONTROL_IN_ACK;
	--			PREV_READ <= PREV_READ XOR RES_EN;
				
	--		END IF;
	--	END IF;
	
	--END PROCESS TO_MCU;
	
	
	--QPE_CONTROL_OUT_TO_MCU(0) <= PREV_ACK;
	--QPE_CONTROL_OUT_TO_MCU(1) <= PREV_READ;

	--State_transitions
	STATE_TRANSITIONS : PROCESS (QPE_CONTROL_IN_CLK,QPE_CONTROL_IN_RSTN)
	BEGIN
	
	IF QPE_CONTROL_IN_RSTN = '0' THEN

		CURRENT_STATE <= RESET;

	ELSE
	
		IF RISING_EDGE(QPE_CONTROL_IN_CLK) THEN
		
			CASE CURRENT_STATE IS
			
				WHEN RESET =>
				
					IF QPE_CONTROL_IN_FROM_MCU(1) = '1' THEN
					
						CURRENT_STATE <= INIT_0_IDLE;
						
					ELSE 
					
						CURRENT_STATE <= RESET;
						
					END IF;
					
				WHEN INIT_0_IDLE =>
				
					IF QPE_CONTROL_IN_FROM_MCU(0) = '1' THEN
						CURRENT_STATE <= INIT_0;
					ELSE
						CURRENT_STATE <= INIT_0_IDLE;
					END IF;
					
					
				WHEN INIT_0 => 
				
					CURRENT_STATE <= INIT_0_END;
					
				WHEN INIT_0_END =>
				
					IF  QPE_CONTROL_IN_FROM_MCU(0) = '0' THEN
						CURRENT_STATE <= INIT_I_IDLE;
					ELSE
						CURRENT_STATE <= INIT_0_END;
					END IF;
					
				WHEN INIT_I_IDLE =>
					
					IF QPE_CONTROL_IN_FROM_MCU(0) = '1' THEN
							CURRENT_STATE <= INIT_I;
					ELSE
							CURRENT_STATE <= INIT_I_IDLE;
					END IF;
		
					
				WHEN INIT_I =>
				
						CURRENT_STATE <= INIT_I_END;
						
				WHEN INIT_I_END =>
					IF  QPE_CONTROL_IN_FROM_MCU(0) = '0' THEN
						CURRENT_STATE <= INIT_II_IDLE;
					ELSE
						CURRENT_STATE <= INIT_I_END;
					END IF;	

					
				
				WHEN INIT_II_IDLE =>
				
					IF QPE_CONTROL_IN_FROM_MCU(1) = '0' THEN
	
						CURRENT_STATE <= START_I_IDLE;

					ELSE 
					
						IF QPE_CONTROL_IN_FROM_MCU(0) = '1' THEN
							CURRENT_STATE <= INIT_II;
						ELSE
							CURRENT_STATE <= INIT_II_IDLE;
						END IF;
						
					END IF;
					
										
				WHEN INIT_II =>
				
						CURRENT_STATE <= INIT_II_END;
				
				WHEN INIT_II_END =>
				
					IF  QPE_CONTROL_IN_FROM_MCU(0) = '0' THEN
						CURRENT_STATE <= INIT_III_IDLE;
					ELSE
						CURRENT_STATE <= INIT_II_END;
					END IF;	
				
				WHEN INIT_III_IDLE =>
					
					IF QPE_CONTROL_IN_FROM_MCU(1) = '0' THEN
	
						CURRENT_STATE <= START_I_IDLE;

					ELSE 
						IF QPE_CONTROL_IN_FROM_MCU(0) = '1' THEN
							CURRENT_STATE <= INIT_III;
						ELSE 
							CURRENT_STATE <= INIT_III_IDLE;
						END IF;
					END IF;		
						
				WHEN INIT_III =>		
					
						CURRENT_STATE <= INIT_III_END;
						
				WHEN INIT_III_END => 
					IF  QPE_CONTROL_IN_FROM_MCU(0) = '0' THEN
						CURRENT_STATE <= INIT_III_IDLE;
					ELSE
						CURRENT_STATE <= INIT_III_END;
					END IF;
					
				WHEN START_I_IDLE =>
					
					IF QPE_CONTROL_IN_FROM_MCU(0) = '1' THEN
						CURRENT_STATE <= START_I;
					ELSE 
						CURRENT_STATE <= START_I_IDLE;
					END IF;
					
					
				WHEN START_I =>
					
					CURRENT_STATE <= START_I_EXE;
					
				WHEN START_I_EXE => 
				
					IF QPE_CONTROL_IN_GATE_COMP = '1' THEN
						CURRENT_STATE <= START_I_END;
					ELSE
						CURRENT_STATE <= START_I_EXE;
					END IF;
				
				WHEN START_I_END =>
				
					IF  QPE_CONTROL_IN_FROM_MCU(0) = '0' THEN
						CURRENT_STATE <= START_II_IDLE;
					ELSE
						CURRENT_STATE <= START_I_END;
					END IF;
				
				WHEN START_II_IDLE =>
				
					IF QPE_CONTROL_IN_FROM_MCU(1) = '1' THEN
	
						CURRENT_STATE <= SEND_IDLE;

					ELSE 
						IF QPE_CONTROL_IN_FROM_MCU(0) = '1' THEN
							CURRENT_STATE <= START_II;
						ELSE 
							CURRENT_STATE <= START_II_IDLE;
						END IF;
					END IF;		
						
				WHEN START_II =>
				
					CURRENT_STATE <= START_II_EXE;
					
				WHEN START_II_EXE =>
				
					IF QPE_CONTROL_IN_GATE_COMP = '1' THEN
						CURRENT_STATE <= START_II_END;
					ELSE
						CURRENT_STATE <= START_II_EXE;
					END IF;
					
				WHEN START_II_END =>
					IF  QPE_CONTROL_IN_FROM_MCU(0) = '0' THEN
						CURRENT_STATE <= START_II_IDLE;
					ELSE
						CURRENT_STATE <= START_II_END;
					END IF;
					
				WHEN SEND_IDLE =>
					
					IF QPE_CONTROL_IN_FROM_MCU(0) = '1' THEN
						CURRENT_STATE <= SEND_END;
					ELSE 
						CURRENT_STATE <= SEND_IDLE;
					END IF;
					
				WHEN SEND =>
				
					CURRENT_STATE <= SEND_IDLE;
					
				WHEN SEND_END =>
				IF QPE_CONTROL_IN_FROM_MCU(0) = '0' THEN
					IF QPE_CONTROL_IN_COMPLETED = '1' THEN
						CURRENT_STATE <= RESET;
					ELSE
						CURRENT_STATE <= SEND;
					END IF;
				ELSE 
					CURRENT_STATE <= SEND_END;
				END IF;
			
				WHEN OTHERS => 
					CURRENT_STATE <= RESET;
								
				END CASE;
		
		END IF;
		
	END IF;
	
	END PROCESS STATE_TRANSITIONS;
	
	--Control generation
	CONTROL_GENERATION : PROCESS (CURRENT_STATE)
	BEGIN
		--Default
		CLR <= '0';
		ACK_INIT <= '0';
		RES_EN <= '0';
		CLR_GATE_COMP <= '0';
		QPE_CONTROL_OUT_CLR_ALL <= '0';
		QPE_CONTROL_OUT_EN_RES_CNT <= '0';
		QPE_CONTROL_OUT_SAMPLE_INSTR <= '0';
		QPE_CONTROL_OUT_SAMPLE_SIN_COS <= '0';
		QPE_CONTROL_OUT_SAVE_QUBIT_NUMB <= '0';
		QPE_CONTROL_OUT_SAVE_SIN_COS <= '0';
		QPE_CONTROL_OUT_EN_QEP_DONE <= '0';
		QPE_CONTROL_OUT_TO_MCU <= "00";
		QPE_CONTROL_OUT_EN_OUT_BUF <= '0';
	
		CASE CURRENT_STATE IS
		
			WHEN RESET =>
				CLR <= '1';
				 CLR_GATE_COMP <= '1';
				QPE_CONTROL_OUT_CLR_ALL <= '1';
				
			WHEN INIT_0 =>
			
			WHEN INIT_0_IDLE =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '1';
				
			WHEN INIT_0_END =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '0';
			
			WHEN INIT_I  =>
				QPE_CONTROL_OUT_SAMPLE_INSTR <= '1';
				QPE_CONTROL_OUT_SAVE_QUBIT_NUMB <= '1';
				
			WHEN INIT_I_IDLE =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '1';
			WHEN INIT_I_END =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '0';
				
			WHEN INIT_II  =>
				QPE_CONTROL_OUT_SAMPLE_SIN_COS <= '1';
				
			WHEN INIT_II_IDLE =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '1';
			WHEN INIT_II_END =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '0';
				
			WHEN INIT_III =>
				QPE_CONTROL_OUT_SAMPLE_SIN_COS <= '1';
				QPE_CONTROL_OUT_SAVE_SIN_COS <= '1';
				
			WHEN INIT_III_IDLE =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '1';
			WHEN INIT_III_END =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '0';
				
			WHEN START_I =>
				QPE_CONTROL_OUT_SAVE_SIN_COS <= '1';
				QPE_CONTROL_OUT_SAMPLE_INSTR <= '1';
				
			WHEN START_I_EXE =>
				QPE_CONTROL_OUT_EN_QEP_DONE <= '1';
				
			WHEN START_I_IDLE =>
				QPE_CONTROL_OUT_TO_MCU(1) <= '1';
				QPE_CONTROL_OUT_TO_MCU(0) <= '1';
			WHEN START_I_END =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '0';
				
			WHEN START_II =>
				--QPE_CONTROL_OUT_EN_QEP_DONE <= '1';
				QPE_CONTROL_OUT_SAMPLE_INSTR <= '1';
				 CLR_GATE_COMP <= '1';
			
			WHEN START_II_EXE =>
				QPE_CONTROL_OUT_EN_QEP_DONE <= '1';
			
			WHEN START_II_IDLE =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '1';
				--QPE_CONTROL_OUT_EN_QEP_DONE <= '1';
			WHEN START_II_END =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '0';
				--QPE_CONTROL_OUT_EN_QEP_DONE <= '1';
			
			WHEN SEND_IDLE =>
				QPE_CONTROL_OUT_TO_MCU(1) <= '1';
				QPE_CONTROL_OUT_TO_MCU(0) <= '0';
				QPE_CONTROL_OUT_EN_OUT_BUF <= '1';
			WHEN SEND_END =>
				QPE_CONTROL_OUT_TO_MCU(0) <= '1';
				QPE_CONTROL_OUT_EN_OUT_BUF <= '1';
			WHEN SEND =>
				QPE_CONTROL_OUT_EN_RES_CNT <= '1';
				QPE_CONTROL_OUT_EN_OUT_BUF <= '1';
				RES_EN <= '1';
		
		
			WHEN OTHERS =>
				CLR <= '1';
				QPE_CONTROL_OUT_CLR_ALL <= '1';
			
		END CASE;
			
			
	
	END PROCESS CONTROL_GENERATION;

END state_machine;
