LIBRARY IEEE;
 USE IEEE.STD_LOGIC_1164.ALL;
 ENTITY state_decoder_N_7 IS
 PORT (
 STATE_DECODER_N_7_IN_QTGT : IN STD_LOGIC_VECTOR( 2 DOWNTO 0);
 STATE_DECODER_N_7_IN_QCTRL : IN STD_LOGIC_VECTOR( 2 DOWNTO 0);
 STATE_DECODER_N_7_IN_OPCODE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
 STATE_DECODER_N_7_IN_SAVE_QBIT_NUMBER : IN STD_LOGIC;
 STATE_DECODER_N_7_IN_CLEAR : IN STD_LOGIC;
 STATE_DECODER_N_7_IN_CLK : IN STD_LOGIC;
 STATE_DECODER_N_7_OUT_MASK_FIRST : OUT STD_LOGIC;  
STATE_DECODER_N_7_OUT_CTRL_MASK : OUT STD_LOGIC_VECTOR ( 127 DOWNTO 0)
 );
 END ENTITY;
ARCHITECTURE generated OF state_decoder_N_7 IS
 COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
SIGNAL TO_SAVE_BUF, FROM_SAVE_BUF : STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL DEC_QCTRL, DEC_USED, QUBIT_USED, QUBIT_MASK, QCTRL_ENABLED_STATES : STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL CLR_SAVE_QUBIT, ctrl_tgt_diff  : STD_LOGIC;
BEGIN
STATE_DECODER_N_7_OUT_MASK_FIRST <= '0' WHEN STATE_DECODER_N_7_IN_OPCODE = "0010" OR STATE_DECODER_N_7_IN_OPCODE = "0100" OR STATE_DECODER_N_7_IN_OPCODE = "0101" OR STATE_DECODER_N_7_IN_OPCODE = "0110" OR STATE_DECODER_N_7_IN_OPCODE = "0111" OR STATE_DECODER_N_7_IN_OPCODE = "1011" ELSE '1';
DEC_QCTRL <= 
"0000001" WHEN STATE_DECODER_N_7_IN_QCTRL = "000" ELSE
"0000010" WHEN STATE_DECODER_N_7_IN_QCTRL = "001" ELSE
"0000100" WHEN STATE_DECODER_N_7_IN_QCTRL = "010" ELSE
"0001000" WHEN STATE_DECODER_N_7_IN_QCTRL = "011" ELSE
"0010000" WHEN STATE_DECODER_N_7_IN_QCTRL = "100" ELSE
"0100000" WHEN STATE_DECODER_N_7_IN_QCTRL = "101" ELSE
"1000000" WHEN STATE_DECODER_N_7_IN_QCTRL = "110" ELSE
(OTHERS => '0');
ctrl_tgt_diff <= '1' WHEN STATE_DECODER_N_7_IN_QCTRL = STATE_DECODER_N_7_IN_QTGT ELSE '0';
QCTRL_ENABLED_STATES <= (OTHERS => '1') WHEN ctrl_tgt_diff = '1' ELSE DEC_QCTRL;
DEC_USED <= 
"0000001" WHEN STATE_DECODER_N_7_IN_QCTRL = "000" ELSE
"0000011" WHEN STATE_DECODER_N_7_IN_QCTRL = "001" ELSE
"0000111" WHEN STATE_DECODER_N_7_IN_QCTRL = "010" ELSE
"0001111" WHEN STATE_DECODER_N_7_IN_QCTRL = "011" ELSE
"0011111" WHEN STATE_DECODER_N_7_IN_QCTRL = "100" ELSE
"0111111" WHEN STATE_DECODER_N_7_IN_QCTRL = "101" ELSE
"1111111" WHEN STATE_DECODER_N_7_IN_QCTRL = "110" ELSE
(OTHERS => '0');
QUBIT_MASK(0) <= QCTRL_ENABLED_STATES(0) ;
QUBIT_MASK(1) <= QCTRL_ENABLED_STATES(1) ;
QUBIT_MASK(2) <= QCTRL_ENABLED_STATES(2) ;
QUBIT_MASK(3) <= QCTRL_ENABLED_STATES(3) ;
QUBIT_MASK(4) <= QCTRL_ENABLED_STATES(4) ;
QUBIT_MASK(5) <= QCTRL_ENABLED_STATES(5) ;
QUBIT_MASK(6) <= QCTRL_ENABLED_STATES(6) ;
TO_SAVE_BUF(0) <= STATE_DECODER_N_7_IN_SAVE_QBIT_NUMBER;
CLR_SAVE_QUBIT <= STATE_DECODER_N_7_IN_CLEAR OR FROM_SAVE_BUF(0);
REG_SAVE_FLAG : n_bit_register
GENERIC MAP (1)
PORT MAP(
												REG_IN_DATA => TO_SAVE_BUF ,
												REG_IN_ENABLE => STATE_DECODER_N_7_IN_SAVE_QBIT_NUMBER ,
												REG_IN_CLEAR => CLR_SAVE_QUBIT ,
												REG_IN_CLK => STATE_DECODER_N_7_IN_CLK ,
												REG_OUT_DATA => FROM_SAVE_BUF);
REG_SAVE_QUBIT_NUMBER : n_bit_register
GENERIC MAP (7)
PORT MAP(
												REG_IN_DATA => DEC_USED ,
												REG_IN_ENABLE => FROM_SAVE_BUF(0) ,
												REG_IN_CLEAR => STATE_DECODER_N_7_IN_CLEAR ,
												REG_IN_CLK => STATE_DECODER_N_7_IN_CLK ,
												REG_OUT_DATA => QUBIT_USED);
STATE_DECODER_N_7_OUT_CTRL_MASK(0) <= ctrl_tgt_diff;
STATE_DECODER_N_7_OUT_CTRL_MASK(1) <= QUBIT_MASK(0);
STATE_DECODER_N_7_OUT_CTRL_MASK(2) <= QUBIT_MASK(1);
STATE_DECODER_N_7_OUT_CTRL_MASK(3) <= QUBIT_MASK(0) OR QUBIT_MASK(1);
STATE_DECODER_N_7_OUT_CTRL_MASK(4) <= QUBIT_MASK(2);
STATE_DECODER_N_7_OUT_CTRL_MASK(5) <= QUBIT_MASK(0) OR QUBIT_MASK(2);
STATE_DECODER_N_7_OUT_CTRL_MASK(6) <= QUBIT_MASK(1) OR QUBIT_MASK(2);
STATE_DECODER_N_7_OUT_CTRL_MASK(7) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2);
STATE_DECODER_N_7_OUT_CTRL_MASK(8) <= QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(9) <= QUBIT_MASK(0) OR QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(10) <= QUBIT_MASK(1) OR QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(11) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(12) <= QUBIT_MASK(2) OR QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(13) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(14) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(15) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3);
STATE_DECODER_N_7_OUT_CTRL_MASK(16) <= QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(17) <= QUBIT_MASK(0) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(18) <= QUBIT_MASK(1) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(19) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(20) <= QUBIT_MASK(2) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(21) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(22) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(23) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(24) <= QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(25) <= QUBIT_MASK(0) OR QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(26) <= QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(27) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(28) <= QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(29) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(30) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(31) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4);
STATE_DECODER_N_7_OUT_CTRL_MASK(32) <= QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(33) <= QUBIT_MASK(0) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(34) <= QUBIT_MASK(1) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(35) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(36) <= QUBIT_MASK(2) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(37) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(38) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(39) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(40) <= QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(41) <= QUBIT_MASK(0) OR QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(42) <= QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(43) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(44) <= QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(45) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(46) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(47) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(48) <= QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(49) <= QUBIT_MASK(0) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(50) <= QUBIT_MASK(1) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(51) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(52) <= QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(53) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(54) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(55) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(56) <= QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(57) <= QUBIT_MASK(0) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(58) <= QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(59) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(60) <= QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(61) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(62) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(63) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5);
STATE_DECODER_N_7_OUT_CTRL_MASK(64) <= QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(65) <= QUBIT_MASK(0) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(66) <= QUBIT_MASK(1) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(67) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(68) <= QUBIT_MASK(2) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(69) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(70) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(71) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(72) <= QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(73) <= QUBIT_MASK(0) OR QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(74) <= QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(75) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(76) <= QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(77) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(78) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(79) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(80) <= QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(81) <= QUBIT_MASK(0) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(82) <= QUBIT_MASK(1) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(83) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(84) <= QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(85) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(86) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(87) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(88) <= QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(89) <= QUBIT_MASK(0) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(90) <= QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(91) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(92) <= QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(93) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(94) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(95) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(96) <= QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(97) <= QUBIT_MASK(0) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(98) <= QUBIT_MASK(1) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(99) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(100) <= QUBIT_MASK(2) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(101) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(102) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(103) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(104) <= QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(105) <= QUBIT_MASK(0) OR QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(106) <= QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(107) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(108) <= QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(109) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(110) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(111) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(112) <= QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(113) <= QUBIT_MASK(0) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(114) <= QUBIT_MASK(1) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(115) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(116) <= QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(117) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(118) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(119) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(120) <= QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(121) <= QUBIT_MASK(0) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(122) <= QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(123) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(124) <= QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(125) <= QUBIT_MASK(0) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(126) <= QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
STATE_DECODER_N_7_OUT_CTRL_MASK(127) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2) OR QUBIT_MASK(3) OR QUBIT_MASK(4) OR QUBIT_MASK(5) OR QUBIT_MASK(6);
END generated;