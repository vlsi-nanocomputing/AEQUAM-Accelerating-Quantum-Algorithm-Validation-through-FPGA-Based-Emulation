LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY multiplier IS 
	GENERIC (K : INTEGER := 20);
	PORT(
		MULTIPLIER_IN_A : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MULTIPLIER_IN_B : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MULTIPLIER_OUT_RES : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0));
END ENTITY;


