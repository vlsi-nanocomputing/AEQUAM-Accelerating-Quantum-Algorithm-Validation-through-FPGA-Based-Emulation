library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_3_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_3_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_3_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_3_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_3_1_IN_SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		MUX_3_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_3_1 IS

BEGIN

	MUX_3_1_OUT_RES <= 
				MUX_3_1_IN_0 WHEN MUX_3_1_IN_SEL = "00" ELSE
				MUX_3_1_IN_1 WHEN MUX_3_1_IN_SEL = "01" ELSE
				MUX_3_1_IN_2 WHEN MUX_3_1_IN_SEL = "10" ELSE
				(OTHERS => '0');


END behavioral;