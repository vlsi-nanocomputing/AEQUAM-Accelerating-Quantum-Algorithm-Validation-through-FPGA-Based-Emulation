LIBRARY IEEE;
 USE IEEE.STD_LOGIC_1164.ALL;
 ENTITY state_decoder_N_3 IS
 PORT (
 STATE_DECODER_N_3_IN_QTGT : IN STD_LOGIC_VECTOR( 1 DOWNTO 0);
 STATE_DECODER_N_3_IN_QCTRL : IN STD_LOGIC_VECTOR( 1 DOWNTO 0);
 STATE_DECODER_N_3_IN_OPCODE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
 STATE_DECODER_N_3_IN_SAVE_QBIT_NUMBER : IN STD_LOGIC;
 STATE_DECODER_N_3_IN_CLEAR : IN STD_LOGIC;
 STATE_DECODER_N_3_IN_CLK : IN STD_LOGIC;
 STATE_DECODER_N_3_OUT_MASK_FIRST : OUT STD_LOGIC;  
STATE_DECODER_N_3_OUT_CTRL_MASK : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0)
 );
 END ENTITY;
ARCHITECTURE generated OF state_decoder_N_3 IS
 COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
SIGNAL TO_SAVE_BUF, FROM_SAVE_BUF : STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL DEC_QCTRL, DEC_USED, QUBIT_USED, QUBIT_MASK, QCTRL_ENABLED_STATES : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL CLR_SAVE_QUBIT, ctrl_tgt_diff  : STD_LOGIC;
BEGIN
STATE_DECODER_N_3_OUT_MASK_FIRST <= '0' WHEN STATE_DECODER_N_3_IN_OPCODE = "0010" OR STATE_DECODER_N_3_IN_OPCODE = "0100" OR STATE_DECODER_N_3_IN_OPCODE = "0101" OR STATE_DECODER_N_3_IN_OPCODE = "0110" OR STATE_DECODER_N_3_IN_OPCODE = "0111" OR STATE_DECODER_N_3_IN_OPCODE = "1011" ELSE '1';
DEC_QCTRL <= 
"001" WHEN STATE_DECODER_N_3_IN_QCTRL = "00" ELSE
"010" WHEN STATE_DECODER_N_3_IN_QCTRL = "01" ELSE
"100" WHEN STATE_DECODER_N_3_IN_QCTRL = "10" ELSE
(OTHERS => '0');
ctrl_tgt_diff <= '1' WHEN STATE_DECODER_N_3_IN_QCTRL = STATE_DECODER_N_3_IN_QTGT ELSE '0';
QCTRL_ENABLED_STATES <= (OTHERS => '1') WHEN ctrl_tgt_diff = '1' ELSE DEC_QCTRL;
DEC_USED <= 
"001" WHEN STATE_DECODER_N_3_IN_QCTRL = "00" ELSE
"011" WHEN STATE_DECODER_N_3_IN_QCTRL = "01" ELSE
"111" WHEN STATE_DECODER_N_3_IN_QCTRL = "10" ELSE
(OTHERS => '0');
QUBIT_MASK(0) <= QCTRL_ENABLED_STATES(0) ;
QUBIT_MASK(1) <= QCTRL_ENABLED_STATES(1) ;
QUBIT_MASK(2) <= QCTRL_ENABLED_STATES(2) ;
TO_SAVE_BUF(0) <= STATE_DECODER_N_3_IN_SAVE_QBIT_NUMBER;
CLR_SAVE_QUBIT <= STATE_DECODER_N_3_IN_CLEAR OR FROM_SAVE_BUF(0);
REG_SAVE_FLAG : n_bit_register
GENERIC MAP (1)
PORT MAP(
												REG_IN_DATA => TO_SAVE_BUF ,
												REG_IN_ENABLE => STATE_DECODER_N_3_IN_SAVE_QBIT_NUMBER ,
												REG_IN_CLEAR => CLR_SAVE_QUBIT ,
												REG_IN_CLK => STATE_DECODER_N_3_IN_CLK ,
												REG_OUT_DATA => FROM_SAVE_BUF);
REG_SAVE_QUBIT_NUMBER : n_bit_register
GENERIC MAP (3)
PORT MAP(
												REG_IN_DATA => DEC_USED ,
												REG_IN_ENABLE => FROM_SAVE_BUF(0) ,
												REG_IN_CLEAR => STATE_DECODER_N_3_IN_CLEAR ,
												REG_IN_CLK => STATE_DECODER_N_3_IN_CLK ,
												REG_OUT_DATA => QUBIT_USED);
STATE_DECODER_N_3_OUT_CTRL_MASK(0) <= ctrl_tgt_diff;
STATE_DECODER_N_3_OUT_CTRL_MASK(1) <= QUBIT_MASK(0);
STATE_DECODER_N_3_OUT_CTRL_MASK(2) <= QUBIT_MASK(1);
STATE_DECODER_N_3_OUT_CTRL_MASK(3) <= QUBIT_MASK(0) OR QUBIT_MASK(1);
STATE_DECODER_N_3_OUT_CTRL_MASK(4) <= QUBIT_MASK(2);
STATE_DECODER_N_3_OUT_CTRL_MASK(5) <= QUBIT_MASK(0) OR QUBIT_MASK(2);
STATE_DECODER_N_3_OUT_CTRL_MASK(6) <= QUBIT_MASK(1) OR QUBIT_MASK(2);
STATE_DECODER_N_3_OUT_CTRL_MASK(7) <= QUBIT_MASK(0) OR QUBIT_MASK(1) OR QUBIT_MASK(2);
END generated;