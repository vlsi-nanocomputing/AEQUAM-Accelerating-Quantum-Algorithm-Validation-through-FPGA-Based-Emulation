library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_1_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_1_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_1_1_IN_SEL : IN STD_LOGIC_VECTOR (-1 DOWNTO 0);
		MUX_1_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_1_1 IS

BEGIN

	MUX_1_1_OUT_RES <= 
				MUX_1_1_IN_0 WHEN MUX_1_1_IN_SEL = "0" ELSE
				(OTHERS => '0');


END behavioral;