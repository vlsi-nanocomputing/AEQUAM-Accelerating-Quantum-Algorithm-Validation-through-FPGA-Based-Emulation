library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY QEP_N_5_W_1_S_0 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		QEP_N_5_W_1_S_0_IN_START : IN STD_LOGIC;
		QEP_N_5_W_1_S_0_IN_QTGT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);  
		QEP_N_5_W_1_S_0_IN_CTRL_MASK : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		QEP_N_5_W_1_S_0_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		QEP_N_5_W_1_S_0_IN_SIN : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_5_W_1_S_0_IN_COS : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_5_W_1_S_0_IN_WIN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		QEP_N_5_W_1_S_0_IN_OUT_STATE_SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		QEP_N_5_W_1_S_0_IN_REAL_IMAG_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		QEP_N_5_W_1_S_0_IN_CLK : IN STD_LOGIC;
		QEP_N_5_W_1_S_0_IN_CLEAR : IN STD_LOGIC;
		QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF : IN STD_LOGIC;
		QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE : IN STD_LOGIC;
		QEP_N_5_W_1_S_0_OUT_DONE : OUT STD_LOGIC;
		QEP_N_5_W_1_S_0_OUT_DATA : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;
ARCHITECTURE generated OF QEP_N_5_W_1_S_0 IS
COMPONENT multiplexer_2_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_2_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		MUX_2_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_5_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_5_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_5_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_5_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_5_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_5_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_5_1_IN_SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		MUX_5_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_32_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_32_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_SEL : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		MUX_32_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register_clear_1 IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT datapath is
    GENERIC (K : INTEGER := 20);	--K represents the chosen parallelism
	PORT(
		--Data signals
		DATAPATH_IN_A : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_B : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_SINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_COSINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_PIPE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_LD : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_MUX_CTRL : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
		DATAPATH_IN_SUB : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		DATAPATH_IN_SAVED : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_CLEAR : IN STD_LOGIC;
		DATAPATH_IN_CLK : IN STD_LOGIC;
		DATAPATH_OUT_A : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_OUT_B : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0));
END COMPONENT;
COMPONENT control_unit IS
 	PORT (
		--Input signals
		CONTROL_UNIT_IN_START : IN STD_LOGIC;
		CONTROL_UNIT_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CONTROL_UNIT_IN_CLK : IN STD_LOGIC;
		CONTROL_UNIT_IN_CLEAR : IN STD_LOGIC;
		CONTROL_UNIT_OUT_PIPE: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_LD : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_MUX_CTRL : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
		CONTROL_UNIT_OUT_SUB : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		CONTROL_UNIT_OUT_SAVED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_DONE : OUT STD_LOGIC);
END COMPONENT;

SIGNAL TO_STATE_REG_0,TO_STATE_REG_1,TO_STATE_REG_2,TO_STATE_REG_3,TO_STATE_REG_4,TO_STATE_REG_5,TO_STATE_REG_6,TO_STATE_REG_7,TO_STATE_REG_8,TO_STATE_REG_9,TO_STATE_REG_10,TO_STATE_REG_11,TO_STATE_REG_12,TO_STATE_REG_13,TO_STATE_REG_14,TO_STATE_REG_15,TO_STATE_REG_16,TO_STATE_REG_17,TO_STATE_REG_18,TO_STATE_REG_19,TO_STATE_REG_20,TO_STATE_REG_21,TO_STATE_REG_22,TO_STATE_REG_23,TO_STATE_REG_24,TO_STATE_REG_25,TO_STATE_REG_26,TO_STATE_REG_27,TO_STATE_REG_28,TO_STATE_REG_29,TO_STATE_REG_30,TO_STATE_REG_31: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_STATE_REG_0,FROM_STATE_REG_1,FROM_STATE_REG_2,FROM_STATE_REG_3,FROM_STATE_REG_4,FROM_STATE_REG_5,FROM_STATE_REG_6,FROM_STATE_REG_7,FROM_STATE_REG_8,FROM_STATE_REG_9,FROM_STATE_REG_10,FROM_STATE_REG_11,FROM_STATE_REG_12,FROM_STATE_REG_13,FROM_STATE_REG_14,FROM_STATE_REG_15,FROM_STATE_REG_16,FROM_STATE_REG_17,FROM_STATE_REG_18,FROM_STATE_REG_19,FROM_STATE_REG_20,FROM_STATE_REG_21,FROM_STATE_REG_22,FROM_STATE_REG_23,FROM_STATE_REG_24,FROM_STATE_REG_25,FROM_STATE_REG_26,FROM_STATE_REG_27,FROM_STATE_REG_28,FROM_STATE_REG_29,FROM_STATE_REG_30,FROM_STATE_REG_31: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_SELECTION_UNIT_0,FROM_SELECTION_UNIT_1,FROM_SELECTION_UNIT_2,FROM_SELECTION_UNIT_3,FROM_SELECTION_UNIT_4,FROM_SELECTION_UNIT_5,FROM_SELECTION_UNIT_6,FROM_SELECTION_UNIT_7,FROM_SELECTION_UNIT_8,FROM_SELECTION_UNIT_9,FROM_SELECTION_UNIT_10,FROM_SELECTION_UNIT_11,FROM_SELECTION_UNIT_12,FROM_SELECTION_UNIT_13,FROM_SELECTION_UNIT_14,FROM_SELECTION_UNIT_15,FROM_SELECTION_UNIT_16,FROM_SELECTION_UNIT_17,FROM_SELECTION_UNIT_18,FROM_SELECTION_UNIT_19,FROM_SELECTION_UNIT_20,FROM_SELECTION_UNIT_21,FROM_SELECTION_UNIT_22,FROM_SELECTION_UNIT_23,FROM_SELECTION_UNIT_24,FROM_SELECTION_UNIT_25,FROM_SELECTION_UNIT_26,FROM_SELECTION_UNIT_27,FROM_SELECTION_UNIT_28,FROM_SELECTION_UNIT_29,FROM_SELECTION_UNIT_30,FROM_SELECTION_UNIT_31: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_0,FROM_WINDOW_1,FROM_WINDOW_2,FROM_WINDOW_3,FROM_WINDOW_4,FROM_WINDOW_5,FROM_WINDOW_6,FROM_WINDOW_7,FROM_WINDOW_8,FROM_WINDOW_9,FROM_WINDOW_10,FROM_WINDOW_11,FROM_WINDOW_12,FROM_WINDOW_13,FROM_WINDOW_14,FROM_WINDOW_15: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL MASKED_INPUT_0,MASKED_INPUT_2,MASKED_INPUT_4,MASKED_INPUT_6,MASKED_INPUT_8,MASKED_INPUT_10,MASKED_INPUT_12,MASKED_INPUT_14: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_DATAPATHS_0,FROM_DATAPATHS_1,FROM_DATAPATHS_2,FROM_DATAPATHS_3,FROM_DATAPATHS_4,FROM_DATAPATHS_5,FROM_DATAPATHS_6,FROM_DATAPATHS_7,FROM_DATAPATHS_8,FROM_DATAPATHS_9,FROM_DATAPATHS_10,FROM_DATAPATHS_11,FROM_DATAPATHS_12,FROM_DATAPATHS_13,FROM_DATAPATHS_14,FROM_DATAPATHS_15: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_CONTROL_UNITS_0,FROM_CONTROL_UNITS_1,FROM_CONTROL_UNITS_2,FROM_CONTROL_UNITS_3,FROM_CONTROL_UNITS_4,FROM_CONTROL_UNITS_5,FROM_CONTROL_UNITS_6,FROM_CONTROL_UNITS_7,FROM_CONTROL_UNITS_8,FROM_CONTROL_UNITS_9,FROM_CONTROL_UNITS_10,FROM_CONTROL_UNITS_11,FROM_CONTROL_UNITS_12,FROM_CONTROL_UNITS_13,FROM_CONTROL_UNITS_14,FROM_CONTROL_UNITS_15: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL UNWINDOWED_0,UNWINDOWED_1,UNWINDOWED_2,UNWINDOWED_3,UNWINDOWED_4,UNWINDOWED_5,UNWINDOWED_6,UNWINDOWED_7,UNWINDOWED_8,UNWINDOWED_9,UNWINDOWED_10,UNWINDOWED_11,UNWINDOWED_12,UNWINDOWED_13,UNWINDOWED_14,UNWINDOWED_15,UNWINDOWED_16,UNWINDOWED_17,UNWINDOWED_18,UNWINDOWED_19,UNWINDOWED_20,UNWINDOWED_21,UNWINDOWED_22,UNWINDOWED_23,UNWINDOWED_24,UNWINDOWED_25,UNWINDOWED_26,UNWINDOWED_27,UNWINDOWED_28,UNWINDOWED_29,UNWINDOWED_30,UNWINDOWED_31: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_DEC_MASK : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL UNWINDOWED_MASK, REORDERED_MASK, STATE_UPDATE_MASK : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL SELECTED_OUTPUT: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_FIRST_CU_DONE : STD_LOGIC;

BEGIN

STATE_REG_0 : n_bit_register_clear_1
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_0 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(0) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_0);
STATE_REG_1 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1);
STATE_REG_2 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_2 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(2) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_2);
STATE_REG_3 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_3 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(3) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_3);
STATE_REG_4 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_4 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(4) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_4);
STATE_REG_5 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_5 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(5) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_5);
STATE_REG_6 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_6 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(6) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_6);
STATE_REG_7 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_7 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(7) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_7);
STATE_REG_8 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_8 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(8) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_8);
STATE_REG_9 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_9 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(9) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_9);
STATE_REG_10 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_10 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(10) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_10);
STATE_REG_11 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_11 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(11) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_11);
STATE_REG_12 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_12 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(12) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_12);
STATE_REG_13 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_13 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(13) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_13);
STATE_REG_14 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_14 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(14) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_14);
STATE_REG_15 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_15 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(15) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_15);
STATE_REG_16 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_16 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(16) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_16);
STATE_REG_17 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_17 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(17) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_17);
STATE_REG_18 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_18 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(18) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_18);
STATE_REG_19 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_19 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(19) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_19);
STATE_REG_20 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_20 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(20) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_20);
STATE_REG_21 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_21 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(21) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_21);
STATE_REG_22 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_22 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(22) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_22);
STATE_REG_23 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_23 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(23) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_23);
STATE_REG_24 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_24 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(24) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_24);
STATE_REG_25 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_25 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(25) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_25);
STATE_REG_26 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_26 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(26) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_26);
STATE_REG_27 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_27 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(27) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_27);
STATE_REG_28 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_28 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(28) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_28);
STATE_REG_29 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_29 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(29) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_29);
STATE_REG_30 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_30 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(30) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_30);
STATE_REG_31 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_31 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(31) ,
												REG_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_31);


MUX_SEL_UNIT_0 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_0 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_0 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_0 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_0 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_0
									);
MUX_SEL_UNIT_1 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_1 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_2 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_4 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_8 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_16 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_1
									);
MUX_SEL_UNIT_2 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_2 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_1 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_1 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_1 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_2
									);
MUX_SEL_UNIT_3 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_3 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_3 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_5 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_9 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_17 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_3
									);
MUX_SEL_UNIT_4 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_4 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_4 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_2 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_2 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_4
									);
MUX_SEL_UNIT_5 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_5 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_6 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_6 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_10 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_18 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_5
									);
MUX_SEL_UNIT_6 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_6 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_5 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_3 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_3 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_6
									);
MUX_SEL_UNIT_7 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_7 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_7 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_7 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_11 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_19 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_7
									);
MUX_SEL_UNIT_8 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_8 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_8 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_8 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_4 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_4 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_8
									);
MUX_SEL_UNIT_9 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_9 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_10 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_12 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_12 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_20 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_9
									);
MUX_SEL_UNIT_10 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_10 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_9 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_9 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_5 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_5 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_10
									);
MUX_SEL_UNIT_11 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_11 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_11 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_13 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_13 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_21 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_11
									);
MUX_SEL_UNIT_12 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_12 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_12 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_10 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_6 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_6 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_12
									);
MUX_SEL_UNIT_13 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_13 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_14 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_14 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_14 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_22 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_13
									);
MUX_SEL_UNIT_14 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_14 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_13 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_11 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_7 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_7 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_14
									);
MUX_SEL_UNIT_15 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_15 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_15 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_15 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_15 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_23 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_15
									);
MUX_SEL_UNIT_16 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_16 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_16 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_16 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_16 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_8 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_16
									);
MUX_SEL_UNIT_17 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_17 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_18 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_20 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_24 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_24 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_17
									);
MUX_SEL_UNIT_18 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_18 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_17 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_17 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_17 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_9 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_18
									);
MUX_SEL_UNIT_19 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_19 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_19 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_21 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_25 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_25 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_19
									);
MUX_SEL_UNIT_20 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_20 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_20 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_18 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_18 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_10 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_20
									);
MUX_SEL_UNIT_21 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_21 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_22 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_22 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_26 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_26 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_21
									);
MUX_SEL_UNIT_22 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_22 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_21 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_19 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_19 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_11 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_22
									);
MUX_SEL_UNIT_23 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_23 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_23 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_23 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_27 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_27 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_23
									);
MUX_SEL_UNIT_24 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_24 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_24 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_24 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_20 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_12 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_24
									);
MUX_SEL_UNIT_25 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_25 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_26 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_28 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_28 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_28 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_25
									);
MUX_SEL_UNIT_26 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_26 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_25 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_25 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_21 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_13 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_26
									);
MUX_SEL_UNIT_27 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_27 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_27 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_29 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_29 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_29 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_27
									);
MUX_SEL_UNIT_28 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_28 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_28 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_26 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_22 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_14 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_28
									);
MUX_SEL_UNIT_29 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_29 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_30 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_30 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_30 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_30 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_29
									);
MUX_SEL_UNIT_30 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_30 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_29 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_27 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_23 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_15 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_30
									);
MUX_SEL_UNIT_31 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => FROM_STATE_REG_31 ,
										MUX_5_1_IN_1 => FROM_STATE_REG_31 ,
										MUX_5_1_IN_2 => FROM_STATE_REG_31 ,
										MUX_5_1_IN_3 => FROM_STATE_REG_31 ,
										MUX_5_1_IN_4 => FROM_STATE_REG_31 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => FROM_SELECTION_UNIT_31
									);

MUX_WINDOWING_UNIT_0 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_0 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_16 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_0
									);
MUX_WINDOWING_UNIT_1 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_1 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_17 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_1
									);
MUX_WINDOWING_UNIT_2 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_2 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_18 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_2
									);
MUX_WINDOWING_UNIT_3 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_3 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_19 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_3
									);
MUX_WINDOWING_UNIT_4 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_4 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_20 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_4
									);
MUX_WINDOWING_UNIT_5 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_5 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_21 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_5
									);
MUX_WINDOWING_UNIT_6 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_6 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_22 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_6
									);
MUX_WINDOWING_UNIT_7 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_7 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_23 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_7
									);
MUX_WINDOWING_UNIT_8 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_8 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_24 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_8
									);
MUX_WINDOWING_UNIT_9 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_9 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_25 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_9
									);
MUX_WINDOWING_UNIT_10 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_10 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_26 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_10
									);
MUX_WINDOWING_UNIT_11 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_11 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_27 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_11
									);
MUX_WINDOWING_UNIT_12 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_12 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_28 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_12
									);
MUX_WINDOWING_UNIT_13 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_13 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_29 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_13
									);
MUX_WINDOWING_UNIT_14 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_14 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_30 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_14
									);
MUX_WINDOWING_UNIT_15 : multiplexer_2_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_2_1_IN_0 => FROM_SELECTION_UNIT_15 ,
										MUX_2_1_IN_1 => FROM_SELECTION_UNIT_31 ,
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_WIN_SEL ,
										MUX_2_1_OUT_RES => FROM_WINDOW_15
									);
MASKED_INPUT_0 <= FROM_WINDOW_0 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_2 <= FROM_WINDOW_2 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_4 <= FROM_WINDOW_4 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_6 <= FROM_WINDOW_6 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_8 <= FROM_WINDOW_8 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_10 <= FROM_WINDOW_10 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_12 <= FROM_WINDOW_12 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_14 <= FROM_WINDOW_14 WHEN QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');

FROM_WINDOW_DEC_MASK <= 
"01" WHEN QEP_N_5_W_1_S_0_IN_WIN_SEL = "0" ELSE
"10" WHEN QEP_N_5_W_1_S_0_IN_WIN_SEL = "1" ELSE
(OTHERS => '0');

UNWINDOWED_MASK(0) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(2) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(3) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(4) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(5) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(6) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(7) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(8) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(9) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(10) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(11) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(12) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(13) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(14) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(15) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(16) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(17) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(18) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(19) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(20) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(21) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(22) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(23) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(24) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(25) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(26) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(27) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(28) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(29) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(30) <= QEP_N_5_W_1_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(31) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(31) <= FROM_WINDOW_DEC_MASK(1);
MUX_REORD_UPDATE_0 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(0 DOWNTO 0) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(0 DOWNTO 0)
									);
MUX_REORD_UPDATE_1 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(2 DOWNTO 2) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(1 DOWNTO 1)
									);
MUX_REORD_UPDATE_2 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(4 DOWNTO 4) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(2 DOWNTO 2)
									);
MUX_REORD_UPDATE_3 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(6 DOWNTO 6) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(3 DOWNTO 3)
									);
MUX_REORD_UPDATE_4 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(8 DOWNTO 8) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(4 DOWNTO 4)
									);
MUX_REORD_UPDATE_5 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(10 DOWNTO 10) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(5 DOWNTO 5)
									);
MUX_REORD_UPDATE_6 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(12 DOWNTO 12) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(6 DOWNTO 6)
									);
MUX_REORD_UPDATE_7 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(14 DOWNTO 14) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(7 DOWNTO 7)
									);
MUX_REORD_UPDATE_8 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(16 DOWNTO 16) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(8 DOWNTO 8)
									);
MUX_REORD_UPDATE_9 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(18 DOWNTO 18) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(9 DOWNTO 9)
									);
MUX_REORD_UPDATE_10 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(20 DOWNTO 20) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(10 DOWNTO 10)
									);
MUX_REORD_UPDATE_11 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(22 DOWNTO 22) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(11 DOWNTO 11)
									);
MUX_REORD_UPDATE_12 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(24 DOWNTO 24) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(12 DOWNTO 12)
									);
MUX_REORD_UPDATE_13 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(26 DOWNTO 26) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(13 DOWNTO 13)
									);
MUX_REORD_UPDATE_14 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(28 DOWNTO 28) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(14 DOWNTO 14)
									);
MUX_REORD_UPDATE_15 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(30 DOWNTO 30) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(15 DOWNTO 15)
									);
MUX_REORD_UPDATE_16 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(1 DOWNTO 1) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(16 DOWNTO 16)
									);
MUX_REORD_UPDATE_17 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(3 DOWNTO 3) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(17 DOWNTO 17)
									);
MUX_REORD_UPDATE_18 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(5 DOWNTO 5) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(18 DOWNTO 18)
									);
MUX_REORD_UPDATE_19 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(7 DOWNTO 7) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(19 DOWNTO 19)
									);
MUX_REORD_UPDATE_20 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(9 DOWNTO 9) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(20 DOWNTO 20)
									);
MUX_REORD_UPDATE_21 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(11 DOWNTO 11) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(21 DOWNTO 21)
									);
MUX_REORD_UPDATE_22 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(13 DOWNTO 13) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(22 DOWNTO 22)
									);
MUX_REORD_UPDATE_23 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(15 DOWNTO 15) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(23 DOWNTO 23)
									);
MUX_REORD_UPDATE_24 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(17 DOWNTO 17) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(24 DOWNTO 24)
									);
MUX_REORD_UPDATE_25 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(19 DOWNTO 19) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(25 DOWNTO 25)
									);
MUX_REORD_UPDATE_26 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(21 DOWNTO 21) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(26 DOWNTO 26)
									);
MUX_REORD_UPDATE_27 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(23 DOWNTO 23) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(27 DOWNTO 27)
									);
MUX_REORD_UPDATE_28 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(25 DOWNTO 25) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(28 DOWNTO 28)
									);
MUX_REORD_UPDATE_29 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(27 DOWNTO 27) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(29 DOWNTO 29)
									);
MUX_REORD_UPDATE_30 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(29 DOWNTO 29) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(30 DOWNTO 30)
									);
MUX_REORD_UPDATE_31 : multiplexer_5_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_5_1_IN_1 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_5_1_IN_2 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_5_1_IN_3 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_5_1_IN_4 => UNWINDOWED_MASK(31 DOWNTO 31) ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => REORDERED_MASK(31 DOWNTO 31)
									);

STATE_UPDATE_MASK(0) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(0) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(0);
STATE_UPDATE_MASK(1) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(1);
STATE_UPDATE_MASK(2) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(2) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(2);
STATE_UPDATE_MASK(3) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(3) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(3);
STATE_UPDATE_MASK(4) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(4) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(4);
STATE_UPDATE_MASK(5) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(5) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(5);
STATE_UPDATE_MASK(6) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(6) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(6);
STATE_UPDATE_MASK(7) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(7) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(7);
STATE_UPDATE_MASK(8) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(8) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(8);
STATE_UPDATE_MASK(9) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(9) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(9);
STATE_UPDATE_MASK(10) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(10) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(10);
STATE_UPDATE_MASK(11) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(11) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(11);
STATE_UPDATE_MASK(12) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(12) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(12);
STATE_UPDATE_MASK(13) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(13) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(13);
STATE_UPDATE_MASK(14) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(14) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(14);
STATE_UPDATE_MASK(15) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(15) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(15);
STATE_UPDATE_MASK(16) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(16) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(16);
STATE_UPDATE_MASK(17) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(17) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(17);
STATE_UPDATE_MASK(18) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(18) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(18);
STATE_UPDATE_MASK(19) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(19) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(19);
STATE_UPDATE_MASK(20) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(20) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(20);
STATE_UPDATE_MASK(21) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(21) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(21);
STATE_UPDATE_MASK(22) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(22) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(22);
STATE_UPDATE_MASK(23) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(23) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(23);
STATE_UPDATE_MASK(24) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(24) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(24);
STATE_UPDATE_MASK(25) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(25) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(25);
STATE_UPDATE_MASK(26) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(26) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(26);
STATE_UPDATE_MASK(27) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(27) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(27);
STATE_UPDATE_MASK(28) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(28) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(28);
STATE_UPDATE_MASK(29) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(29) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(29);
STATE_UPDATE_MASK(30) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(30) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(30);
STATE_UPDATE_MASK(31) <= QEP_N_5_W_1_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(31) AND QEP_N_5_W_1_S_0_IN_CTRL_MASK(31);

QEP_N_5_W_1_S_0_OUT_DONE <= FROM_FIRST_CU_DONE;
CONTROL_UNIT_0 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
		CONTROL_UNIT_OUT_DONE => FROM_FIRST_CU_DONE );
CONTROL_UNIT_1 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0));
CONTROL_UNIT_2 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0));
CONTROL_UNIT_3 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0));
CONTROL_UNIT_4 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_4(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_4(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_4(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_4(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_4(2 DOWNTO 0));
CONTROL_UNIT_5 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_5(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_5(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_5(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_5(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_5(2 DOWNTO 0));
CONTROL_UNIT_6 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_6(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_6(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_6(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_6(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_6(2 DOWNTO 0));
CONTROL_UNIT_7 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_5_W_1_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_5_W_1_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_7(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_7(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_7(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_7(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_7(2 DOWNTO 0));

DATAPATH_0: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_0 ,
            DATAPATH_IN_B => FROM_WINDOW_1 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_0 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1);
DATAPATH_1: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_2 ,
            DATAPATH_IN_B => FROM_WINDOW_3 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_2 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_3);
DATAPATH_2: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_4 ,
            DATAPATH_IN_B => FROM_WINDOW_5 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_4 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_5);
DATAPATH_3: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_6 ,
            DATAPATH_IN_B => FROM_WINDOW_7 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_6 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_7);
DATAPATH_4: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_8 ,
            DATAPATH_IN_B => FROM_WINDOW_9 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_4(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_4(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_4(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_4(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_4(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_8 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_9);
DATAPATH_5: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_10 ,
            DATAPATH_IN_B => FROM_WINDOW_11 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_5(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_5(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_5(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_5(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_5(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_10 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_11);
DATAPATH_6: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_12 ,
            DATAPATH_IN_B => FROM_WINDOW_13 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_6(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_6(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_6(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_6(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_6(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_12 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_13);
DATAPATH_7: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_14 ,
            DATAPATH_IN_B => FROM_WINDOW_15 ,
            DATAPATH_IN_SINE => QEP_N_5_W_1_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_5_W_1_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_7(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_7(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_7(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_7(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_7(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_5_W_1_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_5_W_1_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_14 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_15);

UNWINDOWED_0 <= FROM_DATAPATHS_0;
UNWINDOWED_1 <= FROM_DATAPATHS_1;
UNWINDOWED_2 <= FROM_DATAPATHS_2;
UNWINDOWED_3 <= FROM_DATAPATHS_3;
UNWINDOWED_4 <= FROM_DATAPATHS_4;
UNWINDOWED_5 <= FROM_DATAPATHS_5;
UNWINDOWED_6 <= FROM_DATAPATHS_6;
UNWINDOWED_7 <= FROM_DATAPATHS_7;
UNWINDOWED_8 <= FROM_DATAPATHS_8;
UNWINDOWED_9 <= FROM_DATAPATHS_9;
UNWINDOWED_10 <= FROM_DATAPATHS_10;
UNWINDOWED_11 <= FROM_DATAPATHS_11;
UNWINDOWED_12 <= FROM_DATAPATHS_12;
UNWINDOWED_13 <= FROM_DATAPATHS_13;
UNWINDOWED_14 <= FROM_DATAPATHS_14;
UNWINDOWED_15 <= FROM_DATAPATHS_15;
UNWINDOWED_16 <= FROM_DATAPATHS_0;
UNWINDOWED_17 <= FROM_DATAPATHS_1;
UNWINDOWED_18 <= FROM_DATAPATHS_2;
UNWINDOWED_19 <= FROM_DATAPATHS_3;
UNWINDOWED_20 <= FROM_DATAPATHS_4;
UNWINDOWED_21 <= FROM_DATAPATHS_5;
UNWINDOWED_22 <= FROM_DATAPATHS_6;
UNWINDOWED_23 <= FROM_DATAPATHS_7;
UNWINDOWED_24 <= FROM_DATAPATHS_8;
UNWINDOWED_25 <= FROM_DATAPATHS_9;
UNWINDOWED_26 <= FROM_DATAPATHS_10;
UNWINDOWED_27 <= FROM_DATAPATHS_11;
UNWINDOWED_28 <= FROM_DATAPATHS_12;
UNWINDOWED_29 <= FROM_DATAPATHS_13;
UNWINDOWED_30 <= FROM_DATAPATHS_14;
UNWINDOWED_31 <= FROM_DATAPATHS_15;

MUX_REORD_UNIT_0 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_0 ,
										MUX_5_1_IN_1 => UNWINDOWED_0 ,
										MUX_5_1_IN_2 => UNWINDOWED_0 ,
										MUX_5_1_IN_3 => UNWINDOWED_0 ,
										MUX_5_1_IN_4 => UNWINDOWED_0 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_0
									);
MUX_REORD_UNIT_1 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_1 ,
										MUX_5_1_IN_1 => UNWINDOWED_2 ,
										MUX_5_1_IN_2 => UNWINDOWED_2 ,
										MUX_5_1_IN_3 => UNWINDOWED_2 ,
										MUX_5_1_IN_4 => UNWINDOWED_2 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_1
									);
MUX_REORD_UNIT_2 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_2 ,
										MUX_5_1_IN_1 => UNWINDOWED_1 ,
										MUX_5_1_IN_2 => UNWINDOWED_4 ,
										MUX_5_1_IN_3 => UNWINDOWED_4 ,
										MUX_5_1_IN_4 => UNWINDOWED_4 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_2
									);
MUX_REORD_UNIT_3 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_3 ,
										MUX_5_1_IN_1 => UNWINDOWED_3 ,
										MUX_5_1_IN_2 => UNWINDOWED_6 ,
										MUX_5_1_IN_3 => UNWINDOWED_6 ,
										MUX_5_1_IN_4 => UNWINDOWED_6 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_3
									);
MUX_REORD_UNIT_4 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_4 ,
										MUX_5_1_IN_1 => UNWINDOWED_4 ,
										MUX_5_1_IN_2 => UNWINDOWED_1 ,
										MUX_5_1_IN_3 => UNWINDOWED_8 ,
										MUX_5_1_IN_4 => UNWINDOWED_8 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_4
									);
MUX_REORD_UNIT_5 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_5 ,
										MUX_5_1_IN_1 => UNWINDOWED_6 ,
										MUX_5_1_IN_2 => UNWINDOWED_3 ,
										MUX_5_1_IN_3 => UNWINDOWED_10 ,
										MUX_5_1_IN_4 => UNWINDOWED_10 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_5
									);
MUX_REORD_UNIT_6 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_6 ,
										MUX_5_1_IN_1 => UNWINDOWED_5 ,
										MUX_5_1_IN_2 => UNWINDOWED_5 ,
										MUX_5_1_IN_3 => UNWINDOWED_12 ,
										MUX_5_1_IN_4 => UNWINDOWED_12 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_6
									);
MUX_REORD_UNIT_7 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_7 ,
										MUX_5_1_IN_1 => UNWINDOWED_7 ,
										MUX_5_1_IN_2 => UNWINDOWED_7 ,
										MUX_5_1_IN_3 => UNWINDOWED_14 ,
										MUX_5_1_IN_4 => UNWINDOWED_14 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_7
									);
MUX_REORD_UNIT_8 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_8 ,
										MUX_5_1_IN_1 => UNWINDOWED_8 ,
										MUX_5_1_IN_2 => UNWINDOWED_8 ,
										MUX_5_1_IN_3 => UNWINDOWED_1 ,
										MUX_5_1_IN_4 => UNWINDOWED_16 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_8
									);
MUX_REORD_UNIT_9 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_9 ,
										MUX_5_1_IN_1 => UNWINDOWED_10 ,
										MUX_5_1_IN_2 => UNWINDOWED_10 ,
										MUX_5_1_IN_3 => UNWINDOWED_3 ,
										MUX_5_1_IN_4 => UNWINDOWED_18 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_9
									);
MUX_REORD_UNIT_10 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_10 ,
										MUX_5_1_IN_1 => UNWINDOWED_9 ,
										MUX_5_1_IN_2 => UNWINDOWED_12 ,
										MUX_5_1_IN_3 => UNWINDOWED_5 ,
										MUX_5_1_IN_4 => UNWINDOWED_20 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_10
									);
MUX_REORD_UNIT_11 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_11 ,
										MUX_5_1_IN_1 => UNWINDOWED_11 ,
										MUX_5_1_IN_2 => UNWINDOWED_14 ,
										MUX_5_1_IN_3 => UNWINDOWED_7 ,
										MUX_5_1_IN_4 => UNWINDOWED_22 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_11
									);
MUX_REORD_UNIT_12 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_12 ,
										MUX_5_1_IN_1 => UNWINDOWED_12 ,
										MUX_5_1_IN_2 => UNWINDOWED_9 ,
										MUX_5_1_IN_3 => UNWINDOWED_9 ,
										MUX_5_1_IN_4 => UNWINDOWED_24 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_12
									);
MUX_REORD_UNIT_13 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_13 ,
										MUX_5_1_IN_1 => UNWINDOWED_14 ,
										MUX_5_1_IN_2 => UNWINDOWED_11 ,
										MUX_5_1_IN_3 => UNWINDOWED_11 ,
										MUX_5_1_IN_4 => UNWINDOWED_26 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_13
									);
MUX_REORD_UNIT_14 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_14 ,
										MUX_5_1_IN_1 => UNWINDOWED_13 ,
										MUX_5_1_IN_2 => UNWINDOWED_13 ,
										MUX_5_1_IN_3 => UNWINDOWED_13 ,
										MUX_5_1_IN_4 => UNWINDOWED_28 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_14
									);
MUX_REORD_UNIT_15 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_15 ,
										MUX_5_1_IN_1 => UNWINDOWED_15 ,
										MUX_5_1_IN_2 => UNWINDOWED_15 ,
										MUX_5_1_IN_3 => UNWINDOWED_15 ,
										MUX_5_1_IN_4 => UNWINDOWED_30 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_15
									);
MUX_REORD_UNIT_16 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_16 ,
										MUX_5_1_IN_1 => UNWINDOWED_16 ,
										MUX_5_1_IN_2 => UNWINDOWED_16 ,
										MUX_5_1_IN_3 => UNWINDOWED_16 ,
										MUX_5_1_IN_4 => UNWINDOWED_1 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_16
									);
MUX_REORD_UNIT_17 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_17 ,
										MUX_5_1_IN_1 => UNWINDOWED_18 ,
										MUX_5_1_IN_2 => UNWINDOWED_18 ,
										MUX_5_1_IN_3 => UNWINDOWED_18 ,
										MUX_5_1_IN_4 => UNWINDOWED_3 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_17
									);
MUX_REORD_UNIT_18 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_18 ,
										MUX_5_1_IN_1 => UNWINDOWED_17 ,
										MUX_5_1_IN_2 => UNWINDOWED_20 ,
										MUX_5_1_IN_3 => UNWINDOWED_20 ,
										MUX_5_1_IN_4 => UNWINDOWED_5 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_18
									);
MUX_REORD_UNIT_19 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_19 ,
										MUX_5_1_IN_1 => UNWINDOWED_19 ,
										MUX_5_1_IN_2 => UNWINDOWED_22 ,
										MUX_5_1_IN_3 => UNWINDOWED_22 ,
										MUX_5_1_IN_4 => UNWINDOWED_7 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_19
									);
MUX_REORD_UNIT_20 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_20 ,
										MUX_5_1_IN_1 => UNWINDOWED_20 ,
										MUX_5_1_IN_2 => UNWINDOWED_17 ,
										MUX_5_1_IN_3 => UNWINDOWED_24 ,
										MUX_5_1_IN_4 => UNWINDOWED_9 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_20
									);
MUX_REORD_UNIT_21 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_21 ,
										MUX_5_1_IN_1 => UNWINDOWED_22 ,
										MUX_5_1_IN_2 => UNWINDOWED_19 ,
										MUX_5_1_IN_3 => UNWINDOWED_26 ,
										MUX_5_1_IN_4 => UNWINDOWED_11 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_21
									);
MUX_REORD_UNIT_22 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_22 ,
										MUX_5_1_IN_1 => UNWINDOWED_21 ,
										MUX_5_1_IN_2 => UNWINDOWED_21 ,
										MUX_5_1_IN_3 => UNWINDOWED_28 ,
										MUX_5_1_IN_4 => UNWINDOWED_13 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_22
									);
MUX_REORD_UNIT_23 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_23 ,
										MUX_5_1_IN_1 => UNWINDOWED_23 ,
										MUX_5_1_IN_2 => UNWINDOWED_23 ,
										MUX_5_1_IN_3 => UNWINDOWED_30 ,
										MUX_5_1_IN_4 => UNWINDOWED_15 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_23
									);
MUX_REORD_UNIT_24 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_24 ,
										MUX_5_1_IN_1 => UNWINDOWED_24 ,
										MUX_5_1_IN_2 => UNWINDOWED_24 ,
										MUX_5_1_IN_3 => UNWINDOWED_17 ,
										MUX_5_1_IN_4 => UNWINDOWED_17 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_24
									);
MUX_REORD_UNIT_25 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_25 ,
										MUX_5_1_IN_1 => UNWINDOWED_26 ,
										MUX_5_1_IN_2 => UNWINDOWED_26 ,
										MUX_5_1_IN_3 => UNWINDOWED_19 ,
										MUX_5_1_IN_4 => UNWINDOWED_19 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_25
									);
MUX_REORD_UNIT_26 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_26 ,
										MUX_5_1_IN_1 => UNWINDOWED_25 ,
										MUX_5_1_IN_2 => UNWINDOWED_28 ,
										MUX_5_1_IN_3 => UNWINDOWED_21 ,
										MUX_5_1_IN_4 => UNWINDOWED_21 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_26
									);
MUX_REORD_UNIT_27 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_27 ,
										MUX_5_1_IN_1 => UNWINDOWED_27 ,
										MUX_5_1_IN_2 => UNWINDOWED_30 ,
										MUX_5_1_IN_3 => UNWINDOWED_23 ,
										MUX_5_1_IN_4 => UNWINDOWED_23 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_27
									);
MUX_REORD_UNIT_28 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_28 ,
										MUX_5_1_IN_1 => UNWINDOWED_28 ,
										MUX_5_1_IN_2 => UNWINDOWED_25 ,
										MUX_5_1_IN_3 => UNWINDOWED_25 ,
										MUX_5_1_IN_4 => UNWINDOWED_25 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_28
									);
MUX_REORD_UNIT_29 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_29 ,
										MUX_5_1_IN_1 => UNWINDOWED_30 ,
										MUX_5_1_IN_2 => UNWINDOWED_27 ,
										MUX_5_1_IN_3 => UNWINDOWED_27 ,
										MUX_5_1_IN_4 => UNWINDOWED_27 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_29
									);
MUX_REORD_UNIT_30 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_30 ,
										MUX_5_1_IN_1 => UNWINDOWED_29 ,
										MUX_5_1_IN_2 => UNWINDOWED_29 ,
										MUX_5_1_IN_3 => UNWINDOWED_29 ,
										MUX_5_1_IN_4 => UNWINDOWED_29 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_30
									);
MUX_REORD_UNIT_31 : multiplexer_5_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_5_1_IN_0 => UNWINDOWED_31 ,
										MUX_5_1_IN_1 => UNWINDOWED_31 ,
										MUX_5_1_IN_2 => UNWINDOWED_31 ,
										MUX_5_1_IN_3 => UNWINDOWED_31 ,
										MUX_5_1_IN_4 => UNWINDOWED_31 ,
				                    			MUX_5_1_IN_SEL => QEP_N_5_W_1_S_0_IN_QTGT ,
										MUX_5_1_OUT_RES => TO_STATE_REG_31
									);

MUX_OUTPUT_SELECTION : multiplexer_32_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_32_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_32_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_32_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_32_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_32_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_32_1_IN_5 => FROM_STATE_REG_5 ,
										MUX_32_1_IN_6 => FROM_STATE_REG_6 ,
										MUX_32_1_IN_7 => FROM_STATE_REG_7 ,
										MUX_32_1_IN_8 => FROM_STATE_REG_8 ,
										MUX_32_1_IN_9 => FROM_STATE_REG_9 ,
										MUX_32_1_IN_10 => FROM_STATE_REG_10 ,
										MUX_32_1_IN_11 => FROM_STATE_REG_11 ,
										MUX_32_1_IN_12 => FROM_STATE_REG_12 ,
										MUX_32_1_IN_13 => FROM_STATE_REG_13 ,
										MUX_32_1_IN_14 => FROM_STATE_REG_14 ,
										MUX_32_1_IN_15 => FROM_STATE_REG_15 ,
										MUX_32_1_IN_16 => FROM_STATE_REG_16 ,
										MUX_32_1_IN_17 => FROM_STATE_REG_17 ,
										MUX_32_1_IN_18 => FROM_STATE_REG_18 ,
										MUX_32_1_IN_19 => FROM_STATE_REG_19 ,
										MUX_32_1_IN_20 => FROM_STATE_REG_20 ,
										MUX_32_1_IN_21 => FROM_STATE_REG_21 ,
										MUX_32_1_IN_22 => FROM_STATE_REG_22 ,
										MUX_32_1_IN_23 => FROM_STATE_REG_23 ,
										MUX_32_1_IN_24 => FROM_STATE_REG_24 ,
										MUX_32_1_IN_25 => FROM_STATE_REG_25 ,
										MUX_32_1_IN_26 => FROM_STATE_REG_26 ,
										MUX_32_1_IN_27 => FROM_STATE_REG_27 ,
										MUX_32_1_IN_28 => FROM_STATE_REG_28 ,
										MUX_32_1_IN_29 => FROM_STATE_REG_29 ,
										MUX_32_1_IN_30 => FROM_STATE_REG_30 ,
										MUX_32_1_IN_31 => FROM_STATE_REG_31 ,
				                    			MUX_32_1_IN_SEL => QEP_N_5_W_1_S_0_IN_OUT_STATE_SEL ,
										MUX_32_1_OUT_RES => SELECTED_OUTPUT
									);
MUX_REAL_IMAG_SELECTION : multiplexer_2_1 GENERIC MAP (K => K)
									PORT MAP (
										MUX_2_1_IN_0 => SELECTED_OUTPUT((2*K-1) DOWNTO K),
										MUX_2_1_IN_1 => SELECTED_OUTPUT((K-1) DOWNTO 0),
				                    			MUX_2_1_IN_SEL => QEP_N_5_W_1_S_0_IN_REAL_IMAG_SEL ,
										MUX_2_1_OUT_RES => QEP_N_5_W_1_S_0_OUT_DATA
									);

END generated;