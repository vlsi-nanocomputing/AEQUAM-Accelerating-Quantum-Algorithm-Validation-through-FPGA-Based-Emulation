library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY QEP_N_6_W_3_S_0 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		QEP_N_6_W_3_S_0_IN_START : IN STD_LOGIC;
		QEP_N_6_W_3_S_0_IN_QTGT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);  
		QEP_N_6_W_3_S_0_IN_CTRL_MASK : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		QEP_N_6_W_3_S_0_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		QEP_N_6_W_3_S_0_IN_SIN : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_6_W_3_S_0_IN_COS : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_6_W_3_S_0_IN_WIN_SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		QEP_N_6_W_3_S_0_IN_OUT_STATE_SEL : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		QEP_N_6_W_3_S_0_IN_REAL_IMAG_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		QEP_N_6_W_3_S_0_IN_CLK : IN STD_LOGIC;
		QEP_N_6_W_3_S_0_IN_CLEAR : IN STD_LOGIC;
		QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF : IN STD_LOGIC;
		QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE : IN STD_LOGIC;
		QEP_N_6_W_3_S_0_OUT_DONE : OUT STD_LOGIC;
		QEP_N_6_W_3_S_0_OUT_DATA : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;
ARCHITECTURE generated OF QEP_N_6_W_3_S_0 IS
COMPONENT multiplexer_2_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_2_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		MUX_2_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_6_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_6_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_6_1_IN_SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		MUX_6_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_64_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_64_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_32 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_33 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_34 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_35 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_36 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_37 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_38 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_39 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_40 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_41 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_42 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_43 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_44 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_45 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_46 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_47 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_48 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_49 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_50 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_51 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_52 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_53 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_54 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_55 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_56 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_57 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_58 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_59 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_60 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_61 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_62 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_63 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_64_1_IN_SEL : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		MUX_64_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_8_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_8_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		MUX_8_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register_clear_1 IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT datapath is
    GENERIC (K : INTEGER := 20);	--K represents the chosen parallelism
	PORT(
		--Data signals
		DATAPATH_IN_A : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_B : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_SINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_COSINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_PIPE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_LD : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_MUX_CTRL : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
		DATAPATH_IN_SUB : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		DATAPATH_IN_SAVED : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_CLEAR : IN STD_LOGIC;
		DATAPATH_IN_CLK : IN STD_LOGIC;
		DATAPATH_OUT_A : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_OUT_B : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0));
END COMPONENT;
COMPONENT control_unit IS
 	PORT (
		--Input signals
		CONTROL_UNIT_IN_START : IN STD_LOGIC;
		CONTROL_UNIT_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CONTROL_UNIT_IN_CLK : IN STD_LOGIC;
		CONTROL_UNIT_IN_CLEAR : IN STD_LOGIC;
		CONTROL_UNIT_OUT_PIPE: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_LD : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_MUX_CTRL : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
		CONTROL_UNIT_OUT_SUB : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		CONTROL_UNIT_OUT_SAVED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_DONE : OUT STD_LOGIC);
END COMPONENT;

SIGNAL TO_STATE_REG_0,TO_STATE_REG_1,TO_STATE_REG_2,TO_STATE_REG_3,TO_STATE_REG_4,TO_STATE_REG_5,TO_STATE_REG_6,TO_STATE_REG_7,TO_STATE_REG_8,TO_STATE_REG_9,TO_STATE_REG_10,TO_STATE_REG_11,TO_STATE_REG_12,TO_STATE_REG_13,TO_STATE_REG_14,TO_STATE_REG_15,TO_STATE_REG_16,TO_STATE_REG_17,TO_STATE_REG_18,TO_STATE_REG_19,TO_STATE_REG_20,TO_STATE_REG_21,TO_STATE_REG_22,TO_STATE_REG_23,TO_STATE_REG_24,TO_STATE_REG_25,TO_STATE_REG_26,TO_STATE_REG_27,TO_STATE_REG_28,TO_STATE_REG_29,TO_STATE_REG_30,TO_STATE_REG_31,TO_STATE_REG_32,TO_STATE_REG_33,TO_STATE_REG_34,TO_STATE_REG_35,TO_STATE_REG_36,TO_STATE_REG_37,TO_STATE_REG_38,TO_STATE_REG_39,TO_STATE_REG_40,TO_STATE_REG_41,TO_STATE_REG_42,TO_STATE_REG_43,TO_STATE_REG_44,TO_STATE_REG_45,TO_STATE_REG_46,TO_STATE_REG_47,TO_STATE_REG_48,TO_STATE_REG_49,TO_STATE_REG_50,TO_STATE_REG_51,TO_STATE_REG_52,TO_STATE_REG_53,TO_STATE_REG_54,TO_STATE_REG_55,TO_STATE_REG_56,TO_STATE_REG_57,TO_STATE_REG_58,TO_STATE_REG_59,TO_STATE_REG_60,TO_STATE_REG_61,TO_STATE_REG_62,TO_STATE_REG_63: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_STATE_REG_0,FROM_STATE_REG_1,FROM_STATE_REG_2,FROM_STATE_REG_3,FROM_STATE_REG_4,FROM_STATE_REG_5,FROM_STATE_REG_6,FROM_STATE_REG_7,FROM_STATE_REG_8,FROM_STATE_REG_9,FROM_STATE_REG_10,FROM_STATE_REG_11,FROM_STATE_REG_12,FROM_STATE_REG_13,FROM_STATE_REG_14,FROM_STATE_REG_15,FROM_STATE_REG_16,FROM_STATE_REG_17,FROM_STATE_REG_18,FROM_STATE_REG_19,FROM_STATE_REG_20,FROM_STATE_REG_21,FROM_STATE_REG_22,FROM_STATE_REG_23,FROM_STATE_REG_24,FROM_STATE_REG_25,FROM_STATE_REG_26,FROM_STATE_REG_27,FROM_STATE_REG_28,FROM_STATE_REG_29,FROM_STATE_REG_30,FROM_STATE_REG_31,FROM_STATE_REG_32,FROM_STATE_REG_33,FROM_STATE_REG_34,FROM_STATE_REG_35,FROM_STATE_REG_36,FROM_STATE_REG_37,FROM_STATE_REG_38,FROM_STATE_REG_39,FROM_STATE_REG_40,FROM_STATE_REG_41,FROM_STATE_REG_42,FROM_STATE_REG_43,FROM_STATE_REG_44,FROM_STATE_REG_45,FROM_STATE_REG_46,FROM_STATE_REG_47,FROM_STATE_REG_48,FROM_STATE_REG_49,FROM_STATE_REG_50,FROM_STATE_REG_51,FROM_STATE_REG_52,FROM_STATE_REG_53,FROM_STATE_REG_54,FROM_STATE_REG_55,FROM_STATE_REG_56,FROM_STATE_REG_57,FROM_STATE_REG_58,FROM_STATE_REG_59,FROM_STATE_REG_60,FROM_STATE_REG_61,FROM_STATE_REG_62,FROM_STATE_REG_63: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_SELECTION_UNIT_0,FROM_SELECTION_UNIT_1,FROM_SELECTION_UNIT_2,FROM_SELECTION_UNIT_3,FROM_SELECTION_UNIT_4,FROM_SELECTION_UNIT_5,FROM_SELECTION_UNIT_6,FROM_SELECTION_UNIT_7,FROM_SELECTION_UNIT_8,FROM_SELECTION_UNIT_9,FROM_SELECTION_UNIT_10,FROM_SELECTION_UNIT_11,FROM_SELECTION_UNIT_12,FROM_SELECTION_UNIT_13,FROM_SELECTION_UNIT_14,FROM_SELECTION_UNIT_15,FROM_SELECTION_UNIT_16,FROM_SELECTION_UNIT_17,FROM_SELECTION_UNIT_18,FROM_SELECTION_UNIT_19,FROM_SELECTION_UNIT_20,FROM_SELECTION_UNIT_21,FROM_SELECTION_UNIT_22,FROM_SELECTION_UNIT_23,FROM_SELECTION_UNIT_24,FROM_SELECTION_UNIT_25,FROM_SELECTION_UNIT_26,FROM_SELECTION_UNIT_27,FROM_SELECTION_UNIT_28,FROM_SELECTION_UNIT_29,FROM_SELECTION_UNIT_30,FROM_SELECTION_UNIT_31,FROM_SELECTION_UNIT_32,FROM_SELECTION_UNIT_33,FROM_SELECTION_UNIT_34,FROM_SELECTION_UNIT_35,FROM_SELECTION_UNIT_36,FROM_SELECTION_UNIT_37,FROM_SELECTION_UNIT_38,FROM_SELECTION_UNIT_39,FROM_SELECTION_UNIT_40,FROM_SELECTION_UNIT_41,FROM_SELECTION_UNIT_42,FROM_SELECTION_UNIT_43,FROM_SELECTION_UNIT_44,FROM_SELECTION_UNIT_45,FROM_SELECTION_UNIT_46,FROM_SELECTION_UNIT_47,FROM_SELECTION_UNIT_48,FROM_SELECTION_UNIT_49,FROM_SELECTION_UNIT_50,FROM_SELECTION_UNIT_51,FROM_SELECTION_UNIT_52,FROM_SELECTION_UNIT_53,FROM_SELECTION_UNIT_54,FROM_SELECTION_UNIT_55,FROM_SELECTION_UNIT_56,FROM_SELECTION_UNIT_57,FROM_SELECTION_UNIT_58,FROM_SELECTION_UNIT_59,FROM_SELECTION_UNIT_60,FROM_SELECTION_UNIT_61,FROM_SELECTION_UNIT_62,FROM_SELECTION_UNIT_63: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_0,FROM_WINDOW_1,FROM_WINDOW_2,FROM_WINDOW_3,FROM_WINDOW_4,FROM_WINDOW_5,FROM_WINDOW_6,FROM_WINDOW_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL MASKED_INPUT_0,MASKED_INPUT_2,MASKED_INPUT_4,MASKED_INPUT_6: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_DATAPATHS_0,FROM_DATAPATHS_1,FROM_DATAPATHS_2,FROM_DATAPATHS_3,FROM_DATAPATHS_4,FROM_DATAPATHS_5,FROM_DATAPATHS_6,FROM_DATAPATHS_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_CONTROL_UNITS_0,FROM_CONTROL_UNITS_1,FROM_CONTROL_UNITS_2,FROM_CONTROL_UNITS_3,FROM_CONTROL_UNITS_4,FROM_CONTROL_UNITS_5,FROM_CONTROL_UNITS_6,FROM_CONTROL_UNITS_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL UNWINDOWED_0,UNWINDOWED_1,UNWINDOWED_2,UNWINDOWED_3,UNWINDOWED_4,UNWINDOWED_5,UNWINDOWED_6,UNWINDOWED_7,UNWINDOWED_8,UNWINDOWED_9,UNWINDOWED_10,UNWINDOWED_11,UNWINDOWED_12,UNWINDOWED_13,UNWINDOWED_14,UNWINDOWED_15,UNWINDOWED_16,UNWINDOWED_17,UNWINDOWED_18,UNWINDOWED_19,UNWINDOWED_20,UNWINDOWED_21,UNWINDOWED_22,UNWINDOWED_23,UNWINDOWED_24,UNWINDOWED_25,UNWINDOWED_26,UNWINDOWED_27,UNWINDOWED_28,UNWINDOWED_29,UNWINDOWED_30,UNWINDOWED_31,UNWINDOWED_32,UNWINDOWED_33,UNWINDOWED_34,UNWINDOWED_35,UNWINDOWED_36,UNWINDOWED_37,UNWINDOWED_38,UNWINDOWED_39,UNWINDOWED_40,UNWINDOWED_41,UNWINDOWED_42,UNWINDOWED_43,UNWINDOWED_44,UNWINDOWED_45,UNWINDOWED_46,UNWINDOWED_47,UNWINDOWED_48,UNWINDOWED_49,UNWINDOWED_50,UNWINDOWED_51,UNWINDOWED_52,UNWINDOWED_53,UNWINDOWED_54,UNWINDOWED_55,UNWINDOWED_56,UNWINDOWED_57,UNWINDOWED_58,UNWINDOWED_59,UNWINDOWED_60,UNWINDOWED_61,UNWINDOWED_62,UNWINDOWED_63: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_DEC_MASK : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL UNWINDOWED_MASK, REORDERED_MASK, STATE_UPDATE_MASK : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL SELECTED_OUTPUT: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_FIRST_CU_DONE : STD_LOGIC;

BEGIN

STATE_REG_0 : n_bit_register_clear_1
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_0 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(0) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_0);
STATE_REG_1 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1);
STATE_REG_2 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_2 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(2) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_2);
STATE_REG_3 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_3 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(3) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_3);
STATE_REG_4 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_4 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(4) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_4);
STATE_REG_5 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_5 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(5) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_5);
STATE_REG_6 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_6 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(6) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_6);
STATE_REG_7 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_7 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(7) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_7);
STATE_REG_8 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_8 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(8) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_8);
STATE_REG_9 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_9 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(9) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_9);
STATE_REG_10 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_10 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(10) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_10);
STATE_REG_11 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_11 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(11) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_11);
STATE_REG_12 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_12 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(12) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_12);
STATE_REG_13 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_13 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(13) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_13);
STATE_REG_14 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_14 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(14) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_14);
STATE_REG_15 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_15 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(15) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_15);
STATE_REG_16 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_16 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(16) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_16);
STATE_REG_17 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_17 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(17) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_17);
STATE_REG_18 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_18 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(18) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_18);
STATE_REG_19 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_19 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(19) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_19);
STATE_REG_20 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_20 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(20) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_20);
STATE_REG_21 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_21 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(21) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_21);
STATE_REG_22 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_22 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(22) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_22);
STATE_REG_23 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_23 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(23) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_23);
STATE_REG_24 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_24 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(24) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_24);
STATE_REG_25 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_25 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(25) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_25);
STATE_REG_26 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_26 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(26) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_26);
STATE_REG_27 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_27 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(27) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_27);
STATE_REG_28 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_28 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(28) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_28);
STATE_REG_29 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_29 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(29) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_29);
STATE_REG_30 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_30 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(30) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_30);
STATE_REG_31 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_31 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(31) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_31);
STATE_REG_32 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_32 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(32) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_32);
STATE_REG_33 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_33 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(33) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_33);
STATE_REG_34 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_34 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(34) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_34);
STATE_REG_35 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_35 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(35) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_35);
STATE_REG_36 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_36 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(36) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_36);
STATE_REG_37 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_37 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(37) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_37);
STATE_REG_38 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_38 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(38) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_38);
STATE_REG_39 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_39 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(39) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_39);
STATE_REG_40 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_40 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(40) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_40);
STATE_REG_41 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_41 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(41) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_41);
STATE_REG_42 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_42 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(42) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_42);
STATE_REG_43 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_43 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(43) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_43);
STATE_REG_44 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_44 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(44) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_44);
STATE_REG_45 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_45 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(45) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_45);
STATE_REG_46 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_46 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(46) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_46);
STATE_REG_47 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_47 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(47) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_47);
STATE_REG_48 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_48 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(48) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_48);
STATE_REG_49 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_49 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(49) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_49);
STATE_REG_50 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_50 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(50) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_50);
STATE_REG_51 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_51 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(51) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_51);
STATE_REG_52 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_52 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(52) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_52);
STATE_REG_53 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_53 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(53) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_53);
STATE_REG_54 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_54 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(54) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_54);
STATE_REG_55 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_55 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(55) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_55);
STATE_REG_56 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_56 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(56) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_56);
STATE_REG_57 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_57 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(57) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_57);
STATE_REG_58 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_58 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(58) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_58);
STATE_REG_59 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_59 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(59) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_59);
STATE_REG_60 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_60 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(60) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_60);
STATE_REG_61 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_61 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(61) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_61);
STATE_REG_62 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_62 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(62) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_62);
STATE_REG_63 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_63 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(63) ,
												REG_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_63);


MUX_SEL_UNIT_0 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_0 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_0 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_0 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_0 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_0 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_0
									);
MUX_SEL_UNIT_1 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_1 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_2 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_4 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_8 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_16 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_32 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_1
									);
MUX_SEL_UNIT_2 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_2 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_1 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_1 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_1 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_1 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_2
									);
MUX_SEL_UNIT_3 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_3 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_3 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_5 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_9 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_17 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_33 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_3
									);
MUX_SEL_UNIT_4 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_4 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_4 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_2 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_2 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_2 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_4
									);
MUX_SEL_UNIT_5 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_5 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_6 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_6 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_10 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_18 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_34 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_5
									);
MUX_SEL_UNIT_6 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_6 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_5 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_3 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_3 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_3 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_6
									);
MUX_SEL_UNIT_7 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_7 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_7 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_7 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_11 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_19 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_35 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_7
									);
MUX_SEL_UNIT_8 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_8 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_8 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_8 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_4 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_4 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_8
									);
MUX_SEL_UNIT_9 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_9 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_10 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_12 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_12 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_20 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_36 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_9
									);
MUX_SEL_UNIT_10 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_10 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_9 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_9 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_5 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_5 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_5 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_10
									);
MUX_SEL_UNIT_11 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_11 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_11 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_13 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_13 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_21 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_37 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_11
									);
MUX_SEL_UNIT_12 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_12 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_12 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_10 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_6 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_6 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_6 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_12
									);
MUX_SEL_UNIT_13 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_13 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_14 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_14 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_14 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_22 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_38 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_13
									);
MUX_SEL_UNIT_14 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_14 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_13 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_11 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_7 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_7 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_7 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_14
									);
MUX_SEL_UNIT_15 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_15 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_15 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_15 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_15 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_23 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_39 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_15
									);
MUX_SEL_UNIT_16 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_16 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_16 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_16 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_16 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_8 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_8 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_16
									);
MUX_SEL_UNIT_17 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_17 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_18 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_20 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_24 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_24 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_40 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_17
									);
MUX_SEL_UNIT_18 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_18 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_17 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_17 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_17 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_9 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_9 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_18
									);
MUX_SEL_UNIT_19 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_19 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_19 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_21 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_25 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_25 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_41 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_19
									);
MUX_SEL_UNIT_20 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_20 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_20 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_18 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_18 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_10 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_10 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_20
									);
MUX_SEL_UNIT_21 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_21 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_22 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_22 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_26 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_26 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_42 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_21
									);
MUX_SEL_UNIT_22 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_22 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_21 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_19 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_19 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_11 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_11 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_22
									);
MUX_SEL_UNIT_23 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_23 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_23 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_23 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_27 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_27 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_43 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_23
									);
MUX_SEL_UNIT_24 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_24 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_24 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_24 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_20 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_12 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_12 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_24
									);
MUX_SEL_UNIT_25 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_25 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_26 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_28 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_28 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_28 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_44 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_25
									);
MUX_SEL_UNIT_26 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_26 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_25 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_25 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_21 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_13 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_13 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_26
									);
MUX_SEL_UNIT_27 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_27 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_27 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_29 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_29 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_29 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_45 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_27
									);
MUX_SEL_UNIT_28 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_28 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_28 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_26 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_22 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_14 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_14 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_28
									);
MUX_SEL_UNIT_29 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_29 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_30 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_30 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_30 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_30 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_46 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_29
									);
MUX_SEL_UNIT_30 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_30 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_29 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_27 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_23 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_15 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_15 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_30
									);
MUX_SEL_UNIT_31 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_31 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_31 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_31 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_31 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_31 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_47 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_31
									);
MUX_SEL_UNIT_32 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_32 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_32 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_32 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_32 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_32 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_16 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_32
									);
MUX_SEL_UNIT_33 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_33 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_34 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_36 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_40 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_48 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_48 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_33
									);
MUX_SEL_UNIT_34 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_34 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_33 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_33 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_33 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_33 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_17 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_34
									);
MUX_SEL_UNIT_35 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_35 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_35 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_37 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_41 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_49 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_49 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_35
									);
MUX_SEL_UNIT_36 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_36 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_36 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_34 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_34 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_34 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_18 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_36
									);
MUX_SEL_UNIT_37 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_37 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_38 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_38 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_42 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_50 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_50 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_37
									);
MUX_SEL_UNIT_38 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_38 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_37 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_35 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_35 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_35 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_19 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_38
									);
MUX_SEL_UNIT_39 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_39 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_39 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_39 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_43 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_51 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_51 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_39
									);
MUX_SEL_UNIT_40 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_40 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_40 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_40 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_36 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_36 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_20 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_40
									);
MUX_SEL_UNIT_41 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_41 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_42 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_44 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_44 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_52 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_52 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_41
									);
MUX_SEL_UNIT_42 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_42 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_41 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_41 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_37 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_37 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_21 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_42
									);
MUX_SEL_UNIT_43 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_43 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_43 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_45 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_45 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_53 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_53 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_43
									);
MUX_SEL_UNIT_44 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_44 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_44 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_42 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_38 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_38 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_22 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_44
									);
MUX_SEL_UNIT_45 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_45 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_46 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_46 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_46 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_54 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_54 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_45
									);
MUX_SEL_UNIT_46 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_46 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_45 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_43 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_39 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_39 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_23 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_46
									);
MUX_SEL_UNIT_47 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_47 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_47 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_47 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_47 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_55 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_55 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_47
									);
MUX_SEL_UNIT_48 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_48 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_48 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_48 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_48 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_40 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_24 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_48
									);
MUX_SEL_UNIT_49 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_49 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_50 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_52 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_56 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_56 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_56 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_49
									);
MUX_SEL_UNIT_50 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_50 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_49 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_49 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_49 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_41 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_25 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_50
									);
MUX_SEL_UNIT_51 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_51 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_51 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_53 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_57 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_57 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_57 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_51
									);
MUX_SEL_UNIT_52 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_52 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_52 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_50 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_50 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_42 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_26 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_52
									);
MUX_SEL_UNIT_53 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_53 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_54 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_54 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_58 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_58 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_58 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_53
									);
MUX_SEL_UNIT_54 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_54 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_53 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_51 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_51 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_43 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_27 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_54
									);
MUX_SEL_UNIT_55 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_55 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_55 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_55 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_59 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_59 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_59 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_55
									);
MUX_SEL_UNIT_56 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_56 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_56 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_56 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_52 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_44 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_28 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_56
									);
MUX_SEL_UNIT_57 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_57 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_58 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_60 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_60 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_60 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_60 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_57
									);
MUX_SEL_UNIT_58 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_58 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_57 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_57 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_53 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_45 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_29 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_58
									);
MUX_SEL_UNIT_59 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_59 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_59 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_61 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_61 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_61 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_61 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_59
									);
MUX_SEL_UNIT_60 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_60 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_60 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_58 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_54 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_46 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_30 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_60
									);
MUX_SEL_UNIT_61 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_61 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_62 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_62 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_62 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_62 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_62 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_61
									);
MUX_SEL_UNIT_62 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_62 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_61 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_59 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_55 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_47 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_31 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_62
									);
MUX_SEL_UNIT_63 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => FROM_STATE_REG_63 ,
										MUX_6_1_IN_1 => FROM_STATE_REG_63 ,
										MUX_6_1_IN_2 => FROM_STATE_REG_63 ,
										MUX_6_1_IN_3 => FROM_STATE_REG_63 ,
										MUX_6_1_IN_4 => FROM_STATE_REG_63 ,
										MUX_6_1_IN_5 => FROM_STATE_REG_63 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => FROM_SELECTION_UNIT_63
									);

MUX_WINDOWING_UNIT_0 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_0 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_8 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_16 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_24 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_32 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_40 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_48 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_56 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_0
									);
MUX_WINDOWING_UNIT_1 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_1 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_9 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_17 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_25 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_33 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_41 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_49 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_57 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_1
									);
MUX_WINDOWING_UNIT_2 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_2 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_10 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_18 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_26 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_34 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_42 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_50 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_58 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_2
									);
MUX_WINDOWING_UNIT_3 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_3 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_11 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_19 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_27 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_35 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_43 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_51 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_59 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_3
									);
MUX_WINDOWING_UNIT_4 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_4 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_12 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_20 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_28 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_36 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_44 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_52 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_60 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_4
									);
MUX_WINDOWING_UNIT_5 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_5 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_13 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_21 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_29 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_37 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_45 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_53 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_61 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_5
									);
MUX_WINDOWING_UNIT_6 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_6 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_14 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_22 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_30 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_38 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_46 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_54 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_62 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_6
									);
MUX_WINDOWING_UNIT_7 : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_SELECTION_UNIT_7 ,
										MUX_8_1_IN_1 => FROM_SELECTION_UNIT_15 ,
										MUX_8_1_IN_2 => FROM_SELECTION_UNIT_23 ,
										MUX_8_1_IN_3 => FROM_SELECTION_UNIT_31 ,
										MUX_8_1_IN_4 => FROM_SELECTION_UNIT_39 ,
										MUX_8_1_IN_5 => FROM_SELECTION_UNIT_47 ,
										MUX_8_1_IN_6 => FROM_SELECTION_UNIT_55 ,
										MUX_8_1_IN_7 => FROM_SELECTION_UNIT_63 ,
				                    			MUX_8_1_IN_SEL => QEP_N_6_W_3_S_0_IN_WIN_SEL ,
										MUX_8_1_OUT_RES => FROM_WINDOW_7
									);
MASKED_INPUT_0 <= FROM_WINDOW_0 WHEN QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_2 <= FROM_WINDOW_2 WHEN QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_4 <= FROM_WINDOW_4 WHEN QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_6 <= FROM_WINDOW_6 WHEN QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');

FROM_WINDOW_DEC_MASK <= 
"00000001" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "000" ELSE
"00000010" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "001" ELSE
"00000100" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "010" ELSE
"00001000" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "011" ELSE
"00010000" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "100" ELSE
"00100000" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "101" ELSE
"01000000" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "110" ELSE
"10000000" WHEN QEP_N_6_W_3_S_0_IN_WIN_SEL = "111" ELSE
(OTHERS => '0');

UNWINDOWED_MASK(0) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(2) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(3) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(4) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(5) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(6) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(7) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(8) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(9) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(10) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(11) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(12) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(13) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(14) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(15) <= FROM_WINDOW_DEC_MASK(1);
UNWINDOWED_MASK(16) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(17) <= FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(18) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(19) <= FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(20) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(21) <= FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(22) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(23) <= FROM_WINDOW_DEC_MASK(2);
UNWINDOWED_MASK(24) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(25) <= FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(26) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(27) <= FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(28) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(29) <= FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(30) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(31) <= FROM_WINDOW_DEC_MASK(3);
UNWINDOWED_MASK(32) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(33) <= FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(34) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(35) <= FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(36) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(37) <= FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(38) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(39) <= FROM_WINDOW_DEC_MASK(4);
UNWINDOWED_MASK(40) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(41) <= FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(42) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(43) <= FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(44) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(45) <= FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(46) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(47) <= FROM_WINDOW_DEC_MASK(5);
UNWINDOWED_MASK(48) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(49) <= FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(50) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(51) <= FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(52) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(53) <= FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(54) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(55) <= FROM_WINDOW_DEC_MASK(6);
UNWINDOWED_MASK(56) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(57) <= FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(58) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(59) <= FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(60) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(61) <= FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(62) <= QEP_N_6_W_3_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(63) <= FROM_WINDOW_DEC_MASK(7);
UNWINDOWED_MASK(63) <= FROM_WINDOW_DEC_MASK(7);
MUX_REORD_UPDATE_0 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(0 DOWNTO 0) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(0 DOWNTO 0)
									);
MUX_REORD_UPDATE_1 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(2 DOWNTO 2) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(1 DOWNTO 1)
									);
MUX_REORD_UPDATE_2 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(4 DOWNTO 4) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(2 DOWNTO 2)
									);
MUX_REORD_UPDATE_3 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(6 DOWNTO 6) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(3 DOWNTO 3)
									);
MUX_REORD_UPDATE_4 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(8 DOWNTO 8) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(4 DOWNTO 4)
									);
MUX_REORD_UPDATE_5 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(10 DOWNTO 10) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(5 DOWNTO 5)
									);
MUX_REORD_UPDATE_6 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(12 DOWNTO 12) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(6 DOWNTO 6)
									);
MUX_REORD_UPDATE_7 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(14 DOWNTO 14) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(7 DOWNTO 7)
									);
MUX_REORD_UPDATE_8 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(8 DOWNTO 8) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(16 DOWNTO 16) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(8 DOWNTO 8)
									);
MUX_REORD_UPDATE_9 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(18 DOWNTO 18) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(9 DOWNTO 9)
									);
MUX_REORD_UPDATE_10 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(10 DOWNTO 10) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(20 DOWNTO 20) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(10 DOWNTO 10)
									);
MUX_REORD_UPDATE_11 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(22 DOWNTO 22) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(11 DOWNTO 11)
									);
MUX_REORD_UPDATE_12 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(12 DOWNTO 12) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(24 DOWNTO 24) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(12 DOWNTO 12)
									);
MUX_REORD_UPDATE_13 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(26 DOWNTO 26) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(13 DOWNTO 13)
									);
MUX_REORD_UPDATE_14 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(14 DOWNTO 14) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(28 DOWNTO 28) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(14 DOWNTO 14)
									);
MUX_REORD_UPDATE_15 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(30 DOWNTO 30) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(15 DOWNTO 15)
									);
MUX_REORD_UPDATE_16 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(16 DOWNTO 16) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(32 DOWNTO 32) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(16 DOWNTO 16)
									);
MUX_REORD_UPDATE_17 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(34 DOWNTO 34) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(17 DOWNTO 17)
									);
MUX_REORD_UPDATE_18 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(18 DOWNTO 18) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(36 DOWNTO 36) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(18 DOWNTO 18)
									);
MUX_REORD_UPDATE_19 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(38 DOWNTO 38) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(19 DOWNTO 19)
									);
MUX_REORD_UPDATE_20 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(20 DOWNTO 20) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(9 DOWNTO 9) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(40 DOWNTO 40) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(20 DOWNTO 20)
									);
MUX_REORD_UPDATE_21 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(11 DOWNTO 11) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(42 DOWNTO 42) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(21 DOWNTO 21)
									);
MUX_REORD_UPDATE_22 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(22 DOWNTO 22) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(13 DOWNTO 13) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(44 DOWNTO 44) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(22 DOWNTO 22)
									);
MUX_REORD_UPDATE_23 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(15 DOWNTO 15) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(46 DOWNTO 46) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(23 DOWNTO 23)
									);
MUX_REORD_UPDATE_24 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(24 DOWNTO 24) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(17 DOWNTO 17) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(48 DOWNTO 48) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(24 DOWNTO 24)
									);
MUX_REORD_UPDATE_25 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(19 DOWNTO 19) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(50 DOWNTO 50) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(25 DOWNTO 25)
									);
MUX_REORD_UPDATE_26 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(26 DOWNTO 26) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(21 DOWNTO 21) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(52 DOWNTO 52) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(26 DOWNTO 26)
									);
MUX_REORD_UPDATE_27 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(23 DOWNTO 23) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(54 DOWNTO 54) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(27 DOWNTO 27)
									);
MUX_REORD_UPDATE_28 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(28 DOWNTO 28) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(25 DOWNTO 25) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(56 DOWNTO 56) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(28 DOWNTO 28)
									);
MUX_REORD_UPDATE_29 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(27 DOWNTO 27) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(58 DOWNTO 58) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(29 DOWNTO 29)
									);
MUX_REORD_UPDATE_30 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(30 DOWNTO 30) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(29 DOWNTO 29) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(60 DOWNTO 60) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(30 DOWNTO 30)
									);
MUX_REORD_UPDATE_31 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(31 DOWNTO 31) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(62 DOWNTO 62) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(31 DOWNTO 31)
									);
MUX_REORD_UPDATE_32 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(32 DOWNTO 32) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(1 DOWNTO 1) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(32 DOWNTO 32)
									);
MUX_REORD_UPDATE_33 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(3 DOWNTO 3) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(33 DOWNTO 33)
									);
MUX_REORD_UPDATE_34 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(34 DOWNTO 34) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(5 DOWNTO 5) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(34 DOWNTO 34)
									);
MUX_REORD_UPDATE_35 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(7 DOWNTO 7) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(35 DOWNTO 35)
									);
MUX_REORD_UPDATE_36 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(36 DOWNTO 36) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(9 DOWNTO 9) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(36 DOWNTO 36)
									);
MUX_REORD_UPDATE_37 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(11 DOWNTO 11) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(37 DOWNTO 37)
									);
MUX_REORD_UPDATE_38 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(38 DOWNTO 38) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(13 DOWNTO 13) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(38 DOWNTO 38)
									);
MUX_REORD_UPDATE_39 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(15 DOWNTO 15) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(39 DOWNTO 39)
									);
MUX_REORD_UPDATE_40 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(40 DOWNTO 40) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(17 DOWNTO 17) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(40 DOWNTO 40)
									);
MUX_REORD_UPDATE_41 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(19 DOWNTO 19) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(41 DOWNTO 41)
									);
MUX_REORD_UPDATE_42 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(42 DOWNTO 42) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(21 DOWNTO 21) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(42 DOWNTO 42)
									);
MUX_REORD_UPDATE_43 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(23 DOWNTO 23) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(43 DOWNTO 43)
									);
MUX_REORD_UPDATE_44 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(44 DOWNTO 44) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(25 DOWNTO 25) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(44 DOWNTO 44)
									);
MUX_REORD_UPDATE_45 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(27 DOWNTO 27) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(45 DOWNTO 45)
									);
MUX_REORD_UPDATE_46 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(46 DOWNTO 46) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(29 DOWNTO 29) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(46 DOWNTO 46)
									);
MUX_REORD_UPDATE_47 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(31 DOWNTO 31) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(47 DOWNTO 47)
									);
MUX_REORD_UPDATE_48 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(48 DOWNTO 48) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(33 DOWNTO 33) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(33 DOWNTO 33) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(48 DOWNTO 48)
									);
MUX_REORD_UPDATE_49 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(35 DOWNTO 35) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(35 DOWNTO 35) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(49 DOWNTO 49)
									);
MUX_REORD_UPDATE_50 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(50 DOWNTO 50) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(37 DOWNTO 37) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(37 DOWNTO 37) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(50 DOWNTO 50)
									);
MUX_REORD_UPDATE_51 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(39 DOWNTO 39) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(39 DOWNTO 39) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(51 DOWNTO 51)
									);
MUX_REORD_UPDATE_52 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(52 DOWNTO 52) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(41 DOWNTO 41) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(41 DOWNTO 41) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(52 DOWNTO 52)
									);
MUX_REORD_UPDATE_53 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(43 DOWNTO 43) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(43 DOWNTO 43) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(53 DOWNTO 53)
									);
MUX_REORD_UPDATE_54 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(54 DOWNTO 54) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(45 DOWNTO 45) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(45 DOWNTO 45) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(54 DOWNTO 54)
									);
MUX_REORD_UPDATE_55 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(47 DOWNTO 47) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(47 DOWNTO 47) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(55 DOWNTO 55)
									);
MUX_REORD_UPDATE_56 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(56 DOWNTO 56) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(49 DOWNTO 49) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(49 DOWNTO 49) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(56 DOWNTO 56)
									);
MUX_REORD_UPDATE_57 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(51 DOWNTO 51) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(51 DOWNTO 51) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(57 DOWNTO 57)
									);
MUX_REORD_UPDATE_58 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(58 DOWNTO 58) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(53 DOWNTO 53) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(53 DOWNTO 53) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(58 DOWNTO 58)
									);
MUX_REORD_UPDATE_59 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(55 DOWNTO 55) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(55 DOWNTO 55) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(59 DOWNTO 59)
									);
MUX_REORD_UPDATE_60 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(60 DOWNTO 60) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(57 DOWNTO 57) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(57 DOWNTO 57) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(60 DOWNTO 60)
									);
MUX_REORD_UPDATE_61 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(59 DOWNTO 59) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(59 DOWNTO 59) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(61 DOWNTO 61)
									);
MUX_REORD_UPDATE_62 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(62 DOWNTO 62) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(61 DOWNTO 61) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(61 DOWNTO 61) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(62 DOWNTO 62)
									);
MUX_REORD_UPDATE_63 : multiplexer_6_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_6_1_IN_1 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_6_1_IN_2 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_6_1_IN_3 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_6_1_IN_4 => UNWINDOWED_MASK(63 DOWNTO 63) ,
										MUX_6_1_IN_5 => UNWINDOWED_MASK(63 DOWNTO 63) ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => REORDERED_MASK(63 DOWNTO 63)
									);

STATE_UPDATE_MASK(0) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(0) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(0);
STATE_UPDATE_MASK(1) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(1);
STATE_UPDATE_MASK(2) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(2) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(2);
STATE_UPDATE_MASK(3) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(3) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(3);
STATE_UPDATE_MASK(4) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(4) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(4);
STATE_UPDATE_MASK(5) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(5) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(5);
STATE_UPDATE_MASK(6) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(6) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(6);
STATE_UPDATE_MASK(7) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(7) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(7);
STATE_UPDATE_MASK(8) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(8) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(8);
STATE_UPDATE_MASK(9) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(9) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(9);
STATE_UPDATE_MASK(10) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(10) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(10);
STATE_UPDATE_MASK(11) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(11) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(11);
STATE_UPDATE_MASK(12) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(12) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(12);
STATE_UPDATE_MASK(13) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(13) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(13);
STATE_UPDATE_MASK(14) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(14) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(14);
STATE_UPDATE_MASK(15) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(15) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(15);
STATE_UPDATE_MASK(16) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(16) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(16);
STATE_UPDATE_MASK(17) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(17) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(17);
STATE_UPDATE_MASK(18) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(18) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(18);
STATE_UPDATE_MASK(19) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(19) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(19);
STATE_UPDATE_MASK(20) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(20) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(20);
STATE_UPDATE_MASK(21) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(21) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(21);
STATE_UPDATE_MASK(22) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(22) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(22);
STATE_UPDATE_MASK(23) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(23) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(23);
STATE_UPDATE_MASK(24) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(24) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(24);
STATE_UPDATE_MASK(25) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(25) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(25);
STATE_UPDATE_MASK(26) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(26) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(26);
STATE_UPDATE_MASK(27) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(27) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(27);
STATE_UPDATE_MASK(28) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(28) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(28);
STATE_UPDATE_MASK(29) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(29) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(29);
STATE_UPDATE_MASK(30) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(30) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(30);
STATE_UPDATE_MASK(31) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(31) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(31);
STATE_UPDATE_MASK(32) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(32) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(32);
STATE_UPDATE_MASK(33) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(33) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(33);
STATE_UPDATE_MASK(34) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(34) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(34);
STATE_UPDATE_MASK(35) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(35) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(35);
STATE_UPDATE_MASK(36) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(36) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(36);
STATE_UPDATE_MASK(37) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(37) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(37);
STATE_UPDATE_MASK(38) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(38) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(38);
STATE_UPDATE_MASK(39) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(39) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(39);
STATE_UPDATE_MASK(40) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(40) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(40);
STATE_UPDATE_MASK(41) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(41) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(41);
STATE_UPDATE_MASK(42) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(42) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(42);
STATE_UPDATE_MASK(43) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(43) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(43);
STATE_UPDATE_MASK(44) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(44) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(44);
STATE_UPDATE_MASK(45) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(45) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(45);
STATE_UPDATE_MASK(46) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(46) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(46);
STATE_UPDATE_MASK(47) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(47) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(47);
STATE_UPDATE_MASK(48) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(48) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(48);
STATE_UPDATE_MASK(49) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(49) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(49);
STATE_UPDATE_MASK(50) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(50) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(50);
STATE_UPDATE_MASK(51) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(51) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(51);
STATE_UPDATE_MASK(52) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(52) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(52);
STATE_UPDATE_MASK(53) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(53) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(53);
STATE_UPDATE_MASK(54) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(54) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(54);
STATE_UPDATE_MASK(55) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(55) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(55);
STATE_UPDATE_MASK(56) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(56) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(56);
STATE_UPDATE_MASK(57) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(57) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(57);
STATE_UPDATE_MASK(58) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(58) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(58);
STATE_UPDATE_MASK(59) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(59) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(59);
STATE_UPDATE_MASK(60) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(60) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(60);
STATE_UPDATE_MASK(61) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(61) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(61);
STATE_UPDATE_MASK(62) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(62) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(62);
STATE_UPDATE_MASK(63) <= QEP_N_6_W_3_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(63) AND QEP_N_6_W_3_S_0_IN_CTRL_MASK(63);

QEP_N_6_W_3_S_0_OUT_DONE <= FROM_FIRST_CU_DONE;
CONTROL_UNIT_0 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_6_W_3_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_6_W_3_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
		CONTROL_UNIT_OUT_DONE => FROM_FIRST_CU_DONE );
CONTROL_UNIT_1 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_6_W_3_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_6_W_3_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0));
CONTROL_UNIT_2 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_6_W_3_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_6_W_3_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0));
CONTROL_UNIT_3 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_6_W_3_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_6_W_3_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0));

DATAPATH_0: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_0 ,
            DATAPATH_IN_B => FROM_WINDOW_1 ,
            DATAPATH_IN_SINE => QEP_N_6_W_3_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_6_W_3_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_0 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1);
DATAPATH_1: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_2 ,
            DATAPATH_IN_B => FROM_WINDOW_3 ,
            DATAPATH_IN_SINE => QEP_N_6_W_3_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_6_W_3_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_2 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_3);
DATAPATH_2: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_4 ,
            DATAPATH_IN_B => FROM_WINDOW_5 ,
            DATAPATH_IN_SINE => QEP_N_6_W_3_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_6_W_3_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_4 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_5);
DATAPATH_3: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_6 ,
            DATAPATH_IN_B => FROM_WINDOW_7 ,
            DATAPATH_IN_SINE => QEP_N_6_W_3_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_6_W_3_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_6_W_3_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_6_W_3_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_6 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_7);

UNWINDOWED_0 <= FROM_DATAPATHS_0;
UNWINDOWED_1 <= FROM_DATAPATHS_1;
UNWINDOWED_2 <= FROM_DATAPATHS_2;
UNWINDOWED_3 <= FROM_DATAPATHS_3;
UNWINDOWED_4 <= FROM_DATAPATHS_4;
UNWINDOWED_5 <= FROM_DATAPATHS_5;
UNWINDOWED_6 <= FROM_DATAPATHS_6;
UNWINDOWED_7 <= FROM_DATAPATHS_7;
UNWINDOWED_8 <= FROM_DATAPATHS_0;
UNWINDOWED_9 <= FROM_DATAPATHS_1;
UNWINDOWED_10 <= FROM_DATAPATHS_2;
UNWINDOWED_11 <= FROM_DATAPATHS_3;
UNWINDOWED_12 <= FROM_DATAPATHS_4;
UNWINDOWED_13 <= FROM_DATAPATHS_5;
UNWINDOWED_14 <= FROM_DATAPATHS_6;
UNWINDOWED_15 <= FROM_DATAPATHS_7;
UNWINDOWED_16 <= FROM_DATAPATHS_0;
UNWINDOWED_17 <= FROM_DATAPATHS_1;
UNWINDOWED_18 <= FROM_DATAPATHS_2;
UNWINDOWED_19 <= FROM_DATAPATHS_3;
UNWINDOWED_20 <= FROM_DATAPATHS_4;
UNWINDOWED_21 <= FROM_DATAPATHS_5;
UNWINDOWED_22 <= FROM_DATAPATHS_6;
UNWINDOWED_23 <= FROM_DATAPATHS_7;
UNWINDOWED_24 <= FROM_DATAPATHS_0;
UNWINDOWED_25 <= FROM_DATAPATHS_1;
UNWINDOWED_26 <= FROM_DATAPATHS_2;
UNWINDOWED_27 <= FROM_DATAPATHS_3;
UNWINDOWED_28 <= FROM_DATAPATHS_4;
UNWINDOWED_29 <= FROM_DATAPATHS_5;
UNWINDOWED_30 <= FROM_DATAPATHS_6;
UNWINDOWED_31 <= FROM_DATAPATHS_7;
UNWINDOWED_32 <= FROM_DATAPATHS_0;
UNWINDOWED_33 <= FROM_DATAPATHS_1;
UNWINDOWED_34 <= FROM_DATAPATHS_2;
UNWINDOWED_35 <= FROM_DATAPATHS_3;
UNWINDOWED_36 <= FROM_DATAPATHS_4;
UNWINDOWED_37 <= FROM_DATAPATHS_5;
UNWINDOWED_38 <= FROM_DATAPATHS_6;
UNWINDOWED_39 <= FROM_DATAPATHS_7;
UNWINDOWED_40 <= FROM_DATAPATHS_0;
UNWINDOWED_41 <= FROM_DATAPATHS_1;
UNWINDOWED_42 <= FROM_DATAPATHS_2;
UNWINDOWED_43 <= FROM_DATAPATHS_3;
UNWINDOWED_44 <= FROM_DATAPATHS_4;
UNWINDOWED_45 <= FROM_DATAPATHS_5;
UNWINDOWED_46 <= FROM_DATAPATHS_6;
UNWINDOWED_47 <= FROM_DATAPATHS_7;
UNWINDOWED_48 <= FROM_DATAPATHS_0;
UNWINDOWED_49 <= FROM_DATAPATHS_1;
UNWINDOWED_50 <= FROM_DATAPATHS_2;
UNWINDOWED_51 <= FROM_DATAPATHS_3;
UNWINDOWED_52 <= FROM_DATAPATHS_4;
UNWINDOWED_53 <= FROM_DATAPATHS_5;
UNWINDOWED_54 <= FROM_DATAPATHS_6;
UNWINDOWED_55 <= FROM_DATAPATHS_7;
UNWINDOWED_56 <= FROM_DATAPATHS_0;
UNWINDOWED_57 <= FROM_DATAPATHS_1;
UNWINDOWED_58 <= FROM_DATAPATHS_2;
UNWINDOWED_59 <= FROM_DATAPATHS_3;
UNWINDOWED_60 <= FROM_DATAPATHS_4;
UNWINDOWED_61 <= FROM_DATAPATHS_5;
UNWINDOWED_62 <= FROM_DATAPATHS_6;
UNWINDOWED_63 <= FROM_DATAPATHS_7;

MUX_REORD_UNIT_0 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_0 ,
										MUX_6_1_IN_1 => UNWINDOWED_0 ,
										MUX_6_1_IN_2 => UNWINDOWED_0 ,
										MUX_6_1_IN_3 => UNWINDOWED_0 ,
										MUX_6_1_IN_4 => UNWINDOWED_0 ,
										MUX_6_1_IN_5 => UNWINDOWED_0 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_0
									);
MUX_REORD_UNIT_1 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_1 ,
										MUX_6_1_IN_1 => UNWINDOWED_2 ,
										MUX_6_1_IN_2 => UNWINDOWED_2 ,
										MUX_6_1_IN_3 => UNWINDOWED_2 ,
										MUX_6_1_IN_4 => UNWINDOWED_2 ,
										MUX_6_1_IN_5 => UNWINDOWED_2 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_1
									);
MUX_REORD_UNIT_2 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_2 ,
										MUX_6_1_IN_1 => UNWINDOWED_1 ,
										MUX_6_1_IN_2 => UNWINDOWED_4 ,
										MUX_6_1_IN_3 => UNWINDOWED_4 ,
										MUX_6_1_IN_4 => UNWINDOWED_4 ,
										MUX_6_1_IN_5 => UNWINDOWED_4 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_2
									);
MUX_REORD_UNIT_3 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_3 ,
										MUX_6_1_IN_1 => UNWINDOWED_3 ,
										MUX_6_1_IN_2 => UNWINDOWED_6 ,
										MUX_6_1_IN_3 => UNWINDOWED_6 ,
										MUX_6_1_IN_4 => UNWINDOWED_6 ,
										MUX_6_1_IN_5 => UNWINDOWED_6 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_3
									);
MUX_REORD_UNIT_4 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_4 ,
										MUX_6_1_IN_1 => UNWINDOWED_4 ,
										MUX_6_1_IN_2 => UNWINDOWED_1 ,
										MUX_6_1_IN_3 => UNWINDOWED_8 ,
										MUX_6_1_IN_4 => UNWINDOWED_8 ,
										MUX_6_1_IN_5 => UNWINDOWED_8 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_4
									);
MUX_REORD_UNIT_5 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_5 ,
										MUX_6_1_IN_1 => UNWINDOWED_6 ,
										MUX_6_1_IN_2 => UNWINDOWED_3 ,
										MUX_6_1_IN_3 => UNWINDOWED_10 ,
										MUX_6_1_IN_4 => UNWINDOWED_10 ,
										MUX_6_1_IN_5 => UNWINDOWED_10 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_5
									);
MUX_REORD_UNIT_6 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_6 ,
										MUX_6_1_IN_1 => UNWINDOWED_5 ,
										MUX_6_1_IN_2 => UNWINDOWED_5 ,
										MUX_6_1_IN_3 => UNWINDOWED_12 ,
										MUX_6_1_IN_4 => UNWINDOWED_12 ,
										MUX_6_1_IN_5 => UNWINDOWED_12 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_6
									);
MUX_REORD_UNIT_7 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_7 ,
										MUX_6_1_IN_1 => UNWINDOWED_7 ,
										MUX_6_1_IN_2 => UNWINDOWED_7 ,
										MUX_6_1_IN_3 => UNWINDOWED_14 ,
										MUX_6_1_IN_4 => UNWINDOWED_14 ,
										MUX_6_1_IN_5 => UNWINDOWED_14 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_7
									);
MUX_REORD_UNIT_8 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_8 ,
										MUX_6_1_IN_1 => UNWINDOWED_8 ,
										MUX_6_1_IN_2 => UNWINDOWED_8 ,
										MUX_6_1_IN_3 => UNWINDOWED_1 ,
										MUX_6_1_IN_4 => UNWINDOWED_16 ,
										MUX_6_1_IN_5 => UNWINDOWED_16 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_8
									);
MUX_REORD_UNIT_9 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_9 ,
										MUX_6_1_IN_1 => UNWINDOWED_10 ,
										MUX_6_1_IN_2 => UNWINDOWED_10 ,
										MUX_6_1_IN_3 => UNWINDOWED_3 ,
										MUX_6_1_IN_4 => UNWINDOWED_18 ,
										MUX_6_1_IN_5 => UNWINDOWED_18 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_9
									);
MUX_REORD_UNIT_10 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_10 ,
										MUX_6_1_IN_1 => UNWINDOWED_9 ,
										MUX_6_1_IN_2 => UNWINDOWED_12 ,
										MUX_6_1_IN_3 => UNWINDOWED_5 ,
										MUX_6_1_IN_4 => UNWINDOWED_20 ,
										MUX_6_1_IN_5 => UNWINDOWED_20 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_10
									);
MUX_REORD_UNIT_11 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_11 ,
										MUX_6_1_IN_1 => UNWINDOWED_11 ,
										MUX_6_1_IN_2 => UNWINDOWED_14 ,
										MUX_6_1_IN_3 => UNWINDOWED_7 ,
										MUX_6_1_IN_4 => UNWINDOWED_22 ,
										MUX_6_1_IN_5 => UNWINDOWED_22 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_11
									);
MUX_REORD_UNIT_12 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_12 ,
										MUX_6_1_IN_1 => UNWINDOWED_12 ,
										MUX_6_1_IN_2 => UNWINDOWED_9 ,
										MUX_6_1_IN_3 => UNWINDOWED_9 ,
										MUX_6_1_IN_4 => UNWINDOWED_24 ,
										MUX_6_1_IN_5 => UNWINDOWED_24 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_12
									);
MUX_REORD_UNIT_13 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_13 ,
										MUX_6_1_IN_1 => UNWINDOWED_14 ,
										MUX_6_1_IN_2 => UNWINDOWED_11 ,
										MUX_6_1_IN_3 => UNWINDOWED_11 ,
										MUX_6_1_IN_4 => UNWINDOWED_26 ,
										MUX_6_1_IN_5 => UNWINDOWED_26 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_13
									);
MUX_REORD_UNIT_14 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_14 ,
										MUX_6_1_IN_1 => UNWINDOWED_13 ,
										MUX_6_1_IN_2 => UNWINDOWED_13 ,
										MUX_6_1_IN_3 => UNWINDOWED_13 ,
										MUX_6_1_IN_4 => UNWINDOWED_28 ,
										MUX_6_1_IN_5 => UNWINDOWED_28 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_14
									);
MUX_REORD_UNIT_15 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_15 ,
										MUX_6_1_IN_1 => UNWINDOWED_15 ,
										MUX_6_1_IN_2 => UNWINDOWED_15 ,
										MUX_6_1_IN_3 => UNWINDOWED_15 ,
										MUX_6_1_IN_4 => UNWINDOWED_30 ,
										MUX_6_1_IN_5 => UNWINDOWED_30 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_15
									);
MUX_REORD_UNIT_16 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_16 ,
										MUX_6_1_IN_1 => UNWINDOWED_16 ,
										MUX_6_1_IN_2 => UNWINDOWED_16 ,
										MUX_6_1_IN_3 => UNWINDOWED_16 ,
										MUX_6_1_IN_4 => UNWINDOWED_1 ,
										MUX_6_1_IN_5 => UNWINDOWED_32 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_16
									);
MUX_REORD_UNIT_17 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_17 ,
										MUX_6_1_IN_1 => UNWINDOWED_18 ,
										MUX_6_1_IN_2 => UNWINDOWED_18 ,
										MUX_6_1_IN_3 => UNWINDOWED_18 ,
										MUX_6_1_IN_4 => UNWINDOWED_3 ,
										MUX_6_1_IN_5 => UNWINDOWED_34 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_17
									);
MUX_REORD_UNIT_18 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_18 ,
										MUX_6_1_IN_1 => UNWINDOWED_17 ,
										MUX_6_1_IN_2 => UNWINDOWED_20 ,
										MUX_6_1_IN_3 => UNWINDOWED_20 ,
										MUX_6_1_IN_4 => UNWINDOWED_5 ,
										MUX_6_1_IN_5 => UNWINDOWED_36 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_18
									);
MUX_REORD_UNIT_19 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_19 ,
										MUX_6_1_IN_1 => UNWINDOWED_19 ,
										MUX_6_1_IN_2 => UNWINDOWED_22 ,
										MUX_6_1_IN_3 => UNWINDOWED_22 ,
										MUX_6_1_IN_4 => UNWINDOWED_7 ,
										MUX_6_1_IN_5 => UNWINDOWED_38 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_19
									);
MUX_REORD_UNIT_20 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_20 ,
										MUX_6_1_IN_1 => UNWINDOWED_20 ,
										MUX_6_1_IN_2 => UNWINDOWED_17 ,
										MUX_6_1_IN_3 => UNWINDOWED_24 ,
										MUX_6_1_IN_4 => UNWINDOWED_9 ,
										MUX_6_1_IN_5 => UNWINDOWED_40 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_20
									);
MUX_REORD_UNIT_21 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_21 ,
										MUX_6_1_IN_1 => UNWINDOWED_22 ,
										MUX_6_1_IN_2 => UNWINDOWED_19 ,
										MUX_6_1_IN_3 => UNWINDOWED_26 ,
										MUX_6_1_IN_4 => UNWINDOWED_11 ,
										MUX_6_1_IN_5 => UNWINDOWED_42 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_21
									);
MUX_REORD_UNIT_22 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_22 ,
										MUX_6_1_IN_1 => UNWINDOWED_21 ,
										MUX_6_1_IN_2 => UNWINDOWED_21 ,
										MUX_6_1_IN_3 => UNWINDOWED_28 ,
										MUX_6_1_IN_4 => UNWINDOWED_13 ,
										MUX_6_1_IN_5 => UNWINDOWED_44 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_22
									);
MUX_REORD_UNIT_23 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_23 ,
										MUX_6_1_IN_1 => UNWINDOWED_23 ,
										MUX_6_1_IN_2 => UNWINDOWED_23 ,
										MUX_6_1_IN_3 => UNWINDOWED_30 ,
										MUX_6_1_IN_4 => UNWINDOWED_15 ,
										MUX_6_1_IN_5 => UNWINDOWED_46 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_23
									);
MUX_REORD_UNIT_24 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_24 ,
										MUX_6_1_IN_1 => UNWINDOWED_24 ,
										MUX_6_1_IN_2 => UNWINDOWED_24 ,
										MUX_6_1_IN_3 => UNWINDOWED_17 ,
										MUX_6_1_IN_4 => UNWINDOWED_17 ,
										MUX_6_1_IN_5 => UNWINDOWED_48 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_24
									);
MUX_REORD_UNIT_25 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_25 ,
										MUX_6_1_IN_1 => UNWINDOWED_26 ,
										MUX_6_1_IN_2 => UNWINDOWED_26 ,
										MUX_6_1_IN_3 => UNWINDOWED_19 ,
										MUX_6_1_IN_4 => UNWINDOWED_19 ,
										MUX_6_1_IN_5 => UNWINDOWED_50 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_25
									);
MUX_REORD_UNIT_26 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_26 ,
										MUX_6_1_IN_1 => UNWINDOWED_25 ,
										MUX_6_1_IN_2 => UNWINDOWED_28 ,
										MUX_6_1_IN_3 => UNWINDOWED_21 ,
										MUX_6_1_IN_4 => UNWINDOWED_21 ,
										MUX_6_1_IN_5 => UNWINDOWED_52 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_26
									);
MUX_REORD_UNIT_27 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_27 ,
										MUX_6_1_IN_1 => UNWINDOWED_27 ,
										MUX_6_1_IN_2 => UNWINDOWED_30 ,
										MUX_6_1_IN_3 => UNWINDOWED_23 ,
										MUX_6_1_IN_4 => UNWINDOWED_23 ,
										MUX_6_1_IN_5 => UNWINDOWED_54 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_27
									);
MUX_REORD_UNIT_28 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_28 ,
										MUX_6_1_IN_1 => UNWINDOWED_28 ,
										MUX_6_1_IN_2 => UNWINDOWED_25 ,
										MUX_6_1_IN_3 => UNWINDOWED_25 ,
										MUX_6_1_IN_4 => UNWINDOWED_25 ,
										MUX_6_1_IN_5 => UNWINDOWED_56 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_28
									);
MUX_REORD_UNIT_29 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_29 ,
										MUX_6_1_IN_1 => UNWINDOWED_30 ,
										MUX_6_1_IN_2 => UNWINDOWED_27 ,
										MUX_6_1_IN_3 => UNWINDOWED_27 ,
										MUX_6_1_IN_4 => UNWINDOWED_27 ,
										MUX_6_1_IN_5 => UNWINDOWED_58 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_29
									);
MUX_REORD_UNIT_30 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_30 ,
										MUX_6_1_IN_1 => UNWINDOWED_29 ,
										MUX_6_1_IN_2 => UNWINDOWED_29 ,
										MUX_6_1_IN_3 => UNWINDOWED_29 ,
										MUX_6_1_IN_4 => UNWINDOWED_29 ,
										MUX_6_1_IN_5 => UNWINDOWED_60 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_30
									);
MUX_REORD_UNIT_31 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_31 ,
										MUX_6_1_IN_1 => UNWINDOWED_31 ,
										MUX_6_1_IN_2 => UNWINDOWED_31 ,
										MUX_6_1_IN_3 => UNWINDOWED_31 ,
										MUX_6_1_IN_4 => UNWINDOWED_31 ,
										MUX_6_1_IN_5 => UNWINDOWED_62 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_31
									);
MUX_REORD_UNIT_32 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_32 ,
										MUX_6_1_IN_1 => UNWINDOWED_32 ,
										MUX_6_1_IN_2 => UNWINDOWED_32 ,
										MUX_6_1_IN_3 => UNWINDOWED_32 ,
										MUX_6_1_IN_4 => UNWINDOWED_32 ,
										MUX_6_1_IN_5 => UNWINDOWED_1 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_32
									);
MUX_REORD_UNIT_33 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_33 ,
										MUX_6_1_IN_1 => UNWINDOWED_34 ,
										MUX_6_1_IN_2 => UNWINDOWED_34 ,
										MUX_6_1_IN_3 => UNWINDOWED_34 ,
										MUX_6_1_IN_4 => UNWINDOWED_34 ,
										MUX_6_1_IN_5 => UNWINDOWED_3 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_33
									);
MUX_REORD_UNIT_34 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_34 ,
										MUX_6_1_IN_1 => UNWINDOWED_33 ,
										MUX_6_1_IN_2 => UNWINDOWED_36 ,
										MUX_6_1_IN_3 => UNWINDOWED_36 ,
										MUX_6_1_IN_4 => UNWINDOWED_36 ,
										MUX_6_1_IN_5 => UNWINDOWED_5 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_34
									);
MUX_REORD_UNIT_35 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_35 ,
										MUX_6_1_IN_1 => UNWINDOWED_35 ,
										MUX_6_1_IN_2 => UNWINDOWED_38 ,
										MUX_6_1_IN_3 => UNWINDOWED_38 ,
										MUX_6_1_IN_4 => UNWINDOWED_38 ,
										MUX_6_1_IN_5 => UNWINDOWED_7 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_35
									);
MUX_REORD_UNIT_36 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_36 ,
										MUX_6_1_IN_1 => UNWINDOWED_36 ,
										MUX_6_1_IN_2 => UNWINDOWED_33 ,
										MUX_6_1_IN_3 => UNWINDOWED_40 ,
										MUX_6_1_IN_4 => UNWINDOWED_40 ,
										MUX_6_1_IN_5 => UNWINDOWED_9 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_36
									);
MUX_REORD_UNIT_37 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_37 ,
										MUX_6_1_IN_1 => UNWINDOWED_38 ,
										MUX_6_1_IN_2 => UNWINDOWED_35 ,
										MUX_6_1_IN_3 => UNWINDOWED_42 ,
										MUX_6_1_IN_4 => UNWINDOWED_42 ,
										MUX_6_1_IN_5 => UNWINDOWED_11 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_37
									);
MUX_REORD_UNIT_38 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_38 ,
										MUX_6_1_IN_1 => UNWINDOWED_37 ,
										MUX_6_1_IN_2 => UNWINDOWED_37 ,
										MUX_6_1_IN_3 => UNWINDOWED_44 ,
										MUX_6_1_IN_4 => UNWINDOWED_44 ,
										MUX_6_1_IN_5 => UNWINDOWED_13 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_38
									);
MUX_REORD_UNIT_39 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_39 ,
										MUX_6_1_IN_1 => UNWINDOWED_39 ,
										MUX_6_1_IN_2 => UNWINDOWED_39 ,
										MUX_6_1_IN_3 => UNWINDOWED_46 ,
										MUX_6_1_IN_4 => UNWINDOWED_46 ,
										MUX_6_1_IN_5 => UNWINDOWED_15 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_39
									);
MUX_REORD_UNIT_40 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_40 ,
										MUX_6_1_IN_1 => UNWINDOWED_40 ,
										MUX_6_1_IN_2 => UNWINDOWED_40 ,
										MUX_6_1_IN_3 => UNWINDOWED_33 ,
										MUX_6_1_IN_4 => UNWINDOWED_48 ,
										MUX_6_1_IN_5 => UNWINDOWED_17 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_40
									);
MUX_REORD_UNIT_41 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_41 ,
										MUX_6_1_IN_1 => UNWINDOWED_42 ,
										MUX_6_1_IN_2 => UNWINDOWED_42 ,
										MUX_6_1_IN_3 => UNWINDOWED_35 ,
										MUX_6_1_IN_4 => UNWINDOWED_50 ,
										MUX_6_1_IN_5 => UNWINDOWED_19 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_41
									);
MUX_REORD_UNIT_42 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_42 ,
										MUX_6_1_IN_1 => UNWINDOWED_41 ,
										MUX_6_1_IN_2 => UNWINDOWED_44 ,
										MUX_6_1_IN_3 => UNWINDOWED_37 ,
										MUX_6_1_IN_4 => UNWINDOWED_52 ,
										MUX_6_1_IN_5 => UNWINDOWED_21 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_42
									);
MUX_REORD_UNIT_43 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_43 ,
										MUX_6_1_IN_1 => UNWINDOWED_43 ,
										MUX_6_1_IN_2 => UNWINDOWED_46 ,
										MUX_6_1_IN_3 => UNWINDOWED_39 ,
										MUX_6_1_IN_4 => UNWINDOWED_54 ,
										MUX_6_1_IN_5 => UNWINDOWED_23 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_43
									);
MUX_REORD_UNIT_44 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_44 ,
										MUX_6_1_IN_1 => UNWINDOWED_44 ,
										MUX_6_1_IN_2 => UNWINDOWED_41 ,
										MUX_6_1_IN_3 => UNWINDOWED_41 ,
										MUX_6_1_IN_4 => UNWINDOWED_56 ,
										MUX_6_1_IN_5 => UNWINDOWED_25 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_44
									);
MUX_REORD_UNIT_45 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_45 ,
										MUX_6_1_IN_1 => UNWINDOWED_46 ,
										MUX_6_1_IN_2 => UNWINDOWED_43 ,
										MUX_6_1_IN_3 => UNWINDOWED_43 ,
										MUX_6_1_IN_4 => UNWINDOWED_58 ,
										MUX_6_1_IN_5 => UNWINDOWED_27 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_45
									);
MUX_REORD_UNIT_46 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_46 ,
										MUX_6_1_IN_1 => UNWINDOWED_45 ,
										MUX_6_1_IN_2 => UNWINDOWED_45 ,
										MUX_6_1_IN_3 => UNWINDOWED_45 ,
										MUX_6_1_IN_4 => UNWINDOWED_60 ,
										MUX_6_1_IN_5 => UNWINDOWED_29 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_46
									);
MUX_REORD_UNIT_47 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_47 ,
										MUX_6_1_IN_1 => UNWINDOWED_47 ,
										MUX_6_1_IN_2 => UNWINDOWED_47 ,
										MUX_6_1_IN_3 => UNWINDOWED_47 ,
										MUX_6_1_IN_4 => UNWINDOWED_62 ,
										MUX_6_1_IN_5 => UNWINDOWED_31 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_47
									);
MUX_REORD_UNIT_48 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_48 ,
										MUX_6_1_IN_1 => UNWINDOWED_48 ,
										MUX_6_1_IN_2 => UNWINDOWED_48 ,
										MUX_6_1_IN_3 => UNWINDOWED_48 ,
										MUX_6_1_IN_4 => UNWINDOWED_33 ,
										MUX_6_1_IN_5 => UNWINDOWED_33 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_48
									);
MUX_REORD_UNIT_49 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_49 ,
										MUX_6_1_IN_1 => UNWINDOWED_50 ,
										MUX_6_1_IN_2 => UNWINDOWED_50 ,
										MUX_6_1_IN_3 => UNWINDOWED_50 ,
										MUX_6_1_IN_4 => UNWINDOWED_35 ,
										MUX_6_1_IN_5 => UNWINDOWED_35 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_49
									);
MUX_REORD_UNIT_50 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_50 ,
										MUX_6_1_IN_1 => UNWINDOWED_49 ,
										MUX_6_1_IN_2 => UNWINDOWED_52 ,
										MUX_6_1_IN_3 => UNWINDOWED_52 ,
										MUX_6_1_IN_4 => UNWINDOWED_37 ,
										MUX_6_1_IN_5 => UNWINDOWED_37 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_50
									);
MUX_REORD_UNIT_51 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_51 ,
										MUX_6_1_IN_1 => UNWINDOWED_51 ,
										MUX_6_1_IN_2 => UNWINDOWED_54 ,
										MUX_6_1_IN_3 => UNWINDOWED_54 ,
										MUX_6_1_IN_4 => UNWINDOWED_39 ,
										MUX_6_1_IN_5 => UNWINDOWED_39 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_51
									);
MUX_REORD_UNIT_52 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_52 ,
										MUX_6_1_IN_1 => UNWINDOWED_52 ,
										MUX_6_1_IN_2 => UNWINDOWED_49 ,
										MUX_6_1_IN_3 => UNWINDOWED_56 ,
										MUX_6_1_IN_4 => UNWINDOWED_41 ,
										MUX_6_1_IN_5 => UNWINDOWED_41 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_52
									);
MUX_REORD_UNIT_53 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_53 ,
										MUX_6_1_IN_1 => UNWINDOWED_54 ,
										MUX_6_1_IN_2 => UNWINDOWED_51 ,
										MUX_6_1_IN_3 => UNWINDOWED_58 ,
										MUX_6_1_IN_4 => UNWINDOWED_43 ,
										MUX_6_1_IN_5 => UNWINDOWED_43 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_53
									);
MUX_REORD_UNIT_54 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_54 ,
										MUX_6_1_IN_1 => UNWINDOWED_53 ,
										MUX_6_1_IN_2 => UNWINDOWED_53 ,
										MUX_6_1_IN_3 => UNWINDOWED_60 ,
										MUX_6_1_IN_4 => UNWINDOWED_45 ,
										MUX_6_1_IN_5 => UNWINDOWED_45 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_54
									);
MUX_REORD_UNIT_55 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_55 ,
										MUX_6_1_IN_1 => UNWINDOWED_55 ,
										MUX_6_1_IN_2 => UNWINDOWED_55 ,
										MUX_6_1_IN_3 => UNWINDOWED_62 ,
										MUX_6_1_IN_4 => UNWINDOWED_47 ,
										MUX_6_1_IN_5 => UNWINDOWED_47 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_55
									);
MUX_REORD_UNIT_56 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_56 ,
										MUX_6_1_IN_1 => UNWINDOWED_56 ,
										MUX_6_1_IN_2 => UNWINDOWED_56 ,
										MUX_6_1_IN_3 => UNWINDOWED_49 ,
										MUX_6_1_IN_4 => UNWINDOWED_49 ,
										MUX_6_1_IN_5 => UNWINDOWED_49 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_56
									);
MUX_REORD_UNIT_57 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_57 ,
										MUX_6_1_IN_1 => UNWINDOWED_58 ,
										MUX_6_1_IN_2 => UNWINDOWED_58 ,
										MUX_6_1_IN_3 => UNWINDOWED_51 ,
										MUX_6_1_IN_4 => UNWINDOWED_51 ,
										MUX_6_1_IN_5 => UNWINDOWED_51 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_57
									);
MUX_REORD_UNIT_58 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_58 ,
										MUX_6_1_IN_1 => UNWINDOWED_57 ,
										MUX_6_1_IN_2 => UNWINDOWED_60 ,
										MUX_6_1_IN_3 => UNWINDOWED_53 ,
										MUX_6_1_IN_4 => UNWINDOWED_53 ,
										MUX_6_1_IN_5 => UNWINDOWED_53 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_58
									);
MUX_REORD_UNIT_59 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_59 ,
										MUX_6_1_IN_1 => UNWINDOWED_59 ,
										MUX_6_1_IN_2 => UNWINDOWED_62 ,
										MUX_6_1_IN_3 => UNWINDOWED_55 ,
										MUX_6_1_IN_4 => UNWINDOWED_55 ,
										MUX_6_1_IN_5 => UNWINDOWED_55 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_59
									);
MUX_REORD_UNIT_60 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_60 ,
										MUX_6_1_IN_1 => UNWINDOWED_60 ,
										MUX_6_1_IN_2 => UNWINDOWED_57 ,
										MUX_6_1_IN_3 => UNWINDOWED_57 ,
										MUX_6_1_IN_4 => UNWINDOWED_57 ,
										MUX_6_1_IN_5 => UNWINDOWED_57 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_60
									);
MUX_REORD_UNIT_61 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_61 ,
										MUX_6_1_IN_1 => UNWINDOWED_62 ,
										MUX_6_1_IN_2 => UNWINDOWED_59 ,
										MUX_6_1_IN_3 => UNWINDOWED_59 ,
										MUX_6_1_IN_4 => UNWINDOWED_59 ,
										MUX_6_1_IN_5 => UNWINDOWED_59 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_61
									);
MUX_REORD_UNIT_62 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_62 ,
										MUX_6_1_IN_1 => UNWINDOWED_61 ,
										MUX_6_1_IN_2 => UNWINDOWED_61 ,
										MUX_6_1_IN_3 => UNWINDOWED_61 ,
										MUX_6_1_IN_4 => UNWINDOWED_61 ,
										MUX_6_1_IN_5 => UNWINDOWED_61 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_62
									);
MUX_REORD_UNIT_63 : multiplexer_6_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_6_1_IN_0 => UNWINDOWED_63 ,
										MUX_6_1_IN_1 => UNWINDOWED_63 ,
										MUX_6_1_IN_2 => UNWINDOWED_63 ,
										MUX_6_1_IN_3 => UNWINDOWED_63 ,
										MUX_6_1_IN_4 => UNWINDOWED_63 ,
										MUX_6_1_IN_5 => UNWINDOWED_63 ,
				                    			MUX_6_1_IN_SEL => QEP_N_6_W_3_S_0_IN_QTGT ,
										MUX_6_1_OUT_RES => TO_STATE_REG_63
									);

MUX_OUTPUT_SELECTION : multiplexer_64_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_64_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_64_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_64_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_64_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_64_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_64_1_IN_5 => FROM_STATE_REG_5 ,
										MUX_64_1_IN_6 => FROM_STATE_REG_6 ,
										MUX_64_1_IN_7 => FROM_STATE_REG_7 ,
										MUX_64_1_IN_8 => FROM_STATE_REG_8 ,
										MUX_64_1_IN_9 => FROM_STATE_REG_9 ,
										MUX_64_1_IN_10 => FROM_STATE_REG_10 ,
										MUX_64_1_IN_11 => FROM_STATE_REG_11 ,
										MUX_64_1_IN_12 => FROM_STATE_REG_12 ,
										MUX_64_1_IN_13 => FROM_STATE_REG_13 ,
										MUX_64_1_IN_14 => FROM_STATE_REG_14 ,
										MUX_64_1_IN_15 => FROM_STATE_REG_15 ,
										MUX_64_1_IN_16 => FROM_STATE_REG_16 ,
										MUX_64_1_IN_17 => FROM_STATE_REG_17 ,
										MUX_64_1_IN_18 => FROM_STATE_REG_18 ,
										MUX_64_1_IN_19 => FROM_STATE_REG_19 ,
										MUX_64_1_IN_20 => FROM_STATE_REG_20 ,
										MUX_64_1_IN_21 => FROM_STATE_REG_21 ,
										MUX_64_1_IN_22 => FROM_STATE_REG_22 ,
										MUX_64_1_IN_23 => FROM_STATE_REG_23 ,
										MUX_64_1_IN_24 => FROM_STATE_REG_24 ,
										MUX_64_1_IN_25 => FROM_STATE_REG_25 ,
										MUX_64_1_IN_26 => FROM_STATE_REG_26 ,
										MUX_64_1_IN_27 => FROM_STATE_REG_27 ,
										MUX_64_1_IN_28 => FROM_STATE_REG_28 ,
										MUX_64_1_IN_29 => FROM_STATE_REG_29 ,
										MUX_64_1_IN_30 => FROM_STATE_REG_30 ,
										MUX_64_1_IN_31 => FROM_STATE_REG_31 ,
										MUX_64_1_IN_32 => FROM_STATE_REG_32 ,
										MUX_64_1_IN_33 => FROM_STATE_REG_33 ,
										MUX_64_1_IN_34 => FROM_STATE_REG_34 ,
										MUX_64_1_IN_35 => FROM_STATE_REG_35 ,
										MUX_64_1_IN_36 => FROM_STATE_REG_36 ,
										MUX_64_1_IN_37 => FROM_STATE_REG_37 ,
										MUX_64_1_IN_38 => FROM_STATE_REG_38 ,
										MUX_64_1_IN_39 => FROM_STATE_REG_39 ,
										MUX_64_1_IN_40 => FROM_STATE_REG_40 ,
										MUX_64_1_IN_41 => FROM_STATE_REG_41 ,
										MUX_64_1_IN_42 => FROM_STATE_REG_42 ,
										MUX_64_1_IN_43 => FROM_STATE_REG_43 ,
										MUX_64_1_IN_44 => FROM_STATE_REG_44 ,
										MUX_64_1_IN_45 => FROM_STATE_REG_45 ,
										MUX_64_1_IN_46 => FROM_STATE_REG_46 ,
										MUX_64_1_IN_47 => FROM_STATE_REG_47 ,
										MUX_64_1_IN_48 => FROM_STATE_REG_48 ,
										MUX_64_1_IN_49 => FROM_STATE_REG_49 ,
										MUX_64_1_IN_50 => FROM_STATE_REG_50 ,
										MUX_64_1_IN_51 => FROM_STATE_REG_51 ,
										MUX_64_1_IN_52 => FROM_STATE_REG_52 ,
										MUX_64_1_IN_53 => FROM_STATE_REG_53 ,
										MUX_64_1_IN_54 => FROM_STATE_REG_54 ,
										MUX_64_1_IN_55 => FROM_STATE_REG_55 ,
										MUX_64_1_IN_56 => FROM_STATE_REG_56 ,
										MUX_64_1_IN_57 => FROM_STATE_REG_57 ,
										MUX_64_1_IN_58 => FROM_STATE_REG_58 ,
										MUX_64_1_IN_59 => FROM_STATE_REG_59 ,
										MUX_64_1_IN_60 => FROM_STATE_REG_60 ,
										MUX_64_1_IN_61 => FROM_STATE_REG_61 ,
										MUX_64_1_IN_62 => FROM_STATE_REG_62 ,
										MUX_64_1_IN_63 => FROM_STATE_REG_63 ,
				                    			MUX_64_1_IN_SEL => QEP_N_6_W_3_S_0_IN_OUT_STATE_SEL ,
										MUX_64_1_OUT_RES => SELECTED_OUTPUT
									);
MUX_REAL_IMAG_SELECTION : multiplexer_2_1 GENERIC MAP (K => K)
									PORT MAP (
										MUX_2_1_IN_0 => SELECTED_OUTPUT((2*K-1) DOWNTO K),
										MUX_2_1_IN_1 => SELECTED_OUTPUT((K-1) DOWNTO 0),
				                    			MUX_2_1_IN_SEL => QEP_N_6_W_3_S_0_IN_REAL_IMAG_SEL ,
										MUX_2_1_OUT_RES => QEP_N_6_W_3_S_0_OUT_DATA
									);

END generated;