USE WORK.CONTROL_UNIT;

ARCHITECTURE state_machine OF control_unit IS



	--State definition
	TYPE STATE_TYPE IS (IDLE, X_I, Y_I, Z_I, H_I, H_II, H_III, H_IV, S_I, SDG_I, T_I, T_II, T_III, TDG_I, TDG_II, TDG_III, RX_I, RX_II, RX_III, RX_IV, RX_V, RX_VI, RX_VII, RX_VIII, RX_IX, RY_I, RY_II, RY_III, RY_IV, RY_V, RY_VI, RY_VII, RY_VIII, RY_IX, RZ_I, RZ_II, RZ_III, RZ_IV, RZ_V, RZ_VI, RZ_VII, RZ_VIII, RZ_IX, U1_I, U1_II, U1_III, U1_IV, U1_V);
	SIGNAL CURRENT_STATE : STATE_TYPE;

BEGIN 

	--State transition
	STATE_TRANSITION: PROCESS(CONTROL_UNIT_IN_CLK)
	BEGIN
		IF RISING_EDGE(CONTROL_UNIT_IN_CLK) THEN
		
			IF CONTROL_UNIT_IN_CLEAR = '1' THEN
			
				CURRENT_STATE <= IDLE;
			
			ELSE
			
				CASE CURRENT_STATE IS
				
					WHEN 
				
				
				
					WHEN OTHERS => 
									CURRENT_STATE <= IDLE;
				
				END CASE;
			
			END IF;
		
		END IF;
	
	END PROCESS STATE_TRANSITION;

END state_machine;