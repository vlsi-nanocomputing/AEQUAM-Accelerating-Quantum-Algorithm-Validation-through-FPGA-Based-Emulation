LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY non_rot_rom IS 	
	PORT(
		NON_ROT_ROM_IN_ADD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		NON_ROT_ROM_OUT : OUT STD_LOGIC_VECTOR (40 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF non_rot_rom IS

BEGIN

--Output signal follows the pattern
-- |DONE|NEXT_ADD|CTRL_INST|
-- |  1 |  4     |   36    |
--CTRL_INST is divided as follows
-- |PIPE|LD|OBI|OBR|OAI|OAR|S1A|S1B|S2A|S2B|M12A|M1B|M2B|SUB|SAVED|
-- | 3  |3 | 3 | 2 | 2 | 2 | 3 | 2 | 2 | 2 |  1 | 3 | 3 | 2 |  3  |

-- 					   DONE  NEXT_ADD   PIPE    LD      OBI    OBR    OAI    OAR     S1A    S1B    S2A    S2B   M12A    M1B     M2B   SUB     SAVED
-- 						1	     4        3      3       3       2      2      2      3      2 	    2      2     1       3       3     2        3  
	NON_ROT_ROM_OUT <= 
						'1' & "0000" & "000" & "000" & "000" & "11" & "00" & "01" & "000" & "00" & "00" & "00" & '0' & "000" & "000" & "00" & "000"	
						 WHEN NON_ROT_ROM_IN_ADD = "0000" ELSE		--X_I
						
						'1' & "0000" & "000" & "000" & "011" & "01" & "10" & "00" & "000" & "00" & "00" & "00" & '0' & "000" & "000" & "11" & "000"	
						 WHEN NON_ROT_ROM_IN_ADD = "0001" ELSE		--Y_I
						
						'1' & "0000" & "000" & "000" & "001" & "10" & "00" & "00" & "000" & "00" & "00" & "01" & '0' & "000" & "000" & "11" & "000"	
						 WHEN NON_ROT_ROM_IN_ADD = "0010" ELSE		--Z_I
						
						'0' & "1100" & "010" & "000" & "000" & "00" & "00" & "00" & "100" & "00" & "11" & "01" & '0' & "000" & "000" & "00" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "0011" ELSE		--H_I
						
						'1' & "0000" & "000" & "000" & "100" & "01" & "00" & "00" & "000" & "00" & "00" & "01" & '0' & "000" & "000" & "10" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "0100" ELSE		--S_I
						
						'1' & "0000" & "000" & "000" & "010" & "00" & "00" & "00" & "000" & "00" & "00" & "00" & '0' & "000" & "000" & "01" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "0101" ELSE		--SDG_I
						
						'0' & "1000" & "010" & "000" & "000" & "00" & "00" & "00" & "010" & "00" & "10" & "01" & '0' & "000" & "000" & "10" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "0110" ELSE		--T_I
						
						'0' & "1001" & "010" & "000" & "000" & "00" & "00" & "00" & "010" & "00" & "10" & "01" & '0' & "000" & "000" & "01" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "0111" ELSE		--TDG_I
						
						'0' & "1010" & "001" & "000" & "000" & "00" & "00" & "00" & "000" & "00" & "00" & "00" & '1' & "100" & "100" & "00" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "1000" ELSE		--T_II
						
						'0' & "1011" & "001" & "000" & "000" & "00" & "00" & "00" & "000" & "00" & "00" & "00" & '1' & "100" & "100" & "00" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "1001" ELSE		--TDG_II
												
						'1' & "0000" & "000" & "000" & "010" & "01" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "1010" ELSE		--T_III
												
						'1' & "0000" & "000" & "000" & "010" & "01" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "1011" ELSE		--TDG_III
												
						'0' & "1101" & "011" & "000" & "000" & "00" & "00" & "00" & "100" & "00" & "11" & "01" & '1' & "100" & "100" & "11" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "1100" ELSE		--H_II
						
						'0' & "1110" & "001" & "011" & "000" & "00" & "01" & "10" & "001" & "01" & "01" & "10" & '1' & "100" & "100" & "00" & "000"
						 WHEN NON_ROT_ROM_IN_ADD = "1101" ELSE		--H_III
						
						'1' & "0000" & "000" & "000" & "001" & "10" & "00" & "00" & "001" & "01" & "01" & "10" & '0' & "000" & "000" & "00" & "011"
						 WHEN NON_ROT_ROM_IN_ADD = "1110" ELSE		--H_IV
						
						(OTHERS => '0');

END behavioral;