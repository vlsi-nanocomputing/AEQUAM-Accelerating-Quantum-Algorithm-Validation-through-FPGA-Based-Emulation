library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY comb_adder IS 
	GENERIC( K : INTEGER := 20);
	PORT(
		COMB_ADD_IN_A : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		COMB_ADD_IN_B : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		COMB_ADD_IN_CIN : IN STD_LOGIC;
		
		COMB_ADD_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;
