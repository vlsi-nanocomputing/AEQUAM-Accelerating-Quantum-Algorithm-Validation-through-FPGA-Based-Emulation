library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY QEP_N_3_W_0_S_0 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		QEP_N_3_W_0_S_0_IN_START : IN STD_LOGIC;
		QEP_N_3_W_0_S_0_IN_QTGT : IN STD_LOGIC_VECTOR (1 DOWNTO 0);  
		QEP_N_3_W_0_S_0_IN_CTRL_MASK : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		QEP_N_3_W_0_S_0_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		QEP_N_3_W_0_S_0_IN_SIN : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_3_W_0_S_0_IN_COS : IN STD_LOGIC_VECTOR(K-1 DOWNTO 0);
		QEP_N_3_W_0_S_0_IN_OUT_STATE_SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		QEP_N_3_W_0_S_0_IN_REAL_IMAG_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		QEP_N_3_W_0_S_0_IN_CLK : IN STD_LOGIC;
		QEP_N_3_W_0_S_0_IN_CLEAR : IN STD_LOGIC;
		QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF : IN STD_LOGIC;
		QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE : IN STD_LOGIC;
		QEP_N_3_W_0_S_0_OUT_DONE : OUT STD_LOGIC;
		QEP_N_3_W_0_S_0_OUT_DATA : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;
ARCHITECTURE generated OF QEP_N_3_W_0_S_0 IS
COMPONENT multiplexer_2_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_2_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		MUX_2_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_3_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_3_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_3_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_3_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_3_1_IN_SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		MUX_3_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT multiplexer_8_1 IS
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_8_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_8_1_IN_SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		MUX_8_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT n_bit_register_clear_1 IS
	generic (n_bit: INTEGER);
	port (REG_IN_DATA: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    REG_IN_CLK, REG_IN_CLEAR, REG_IN_ENABLE: IN STD_LOGIC;
		    REG_OUT_DATA: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
END COMPONENT;
COMPONENT datapath is
    GENERIC (K : INTEGER := 20);	--K represents the chosen parallelism
	PORT(
		--Data signals
		DATAPATH_IN_A : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_B : IN STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_IN_SINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_COSINE : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		DATAPATH_IN_PIPE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_LD : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_MUX_CTRL : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
		DATAPATH_IN_SUB : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		DATAPATH_IN_SAVED : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DATAPATH_IN_CLEAR : IN STD_LOGIC;
		DATAPATH_IN_CLK : IN STD_LOGIC;
		DATAPATH_OUT_A : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0);
		DATAPATH_OUT_B : OUT STD_LOGIC_VECTOR (2*K-1 DOWNTO 0));
END COMPONENT;
COMPONENT control_unit IS
 	PORT (
		--Input signals
		CONTROL_UNIT_IN_START : IN STD_LOGIC;
		CONTROL_UNIT_IN_OPCODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CONTROL_UNIT_IN_CLK : IN STD_LOGIC;
		CONTROL_UNIT_IN_CLEAR : IN STD_LOGIC;
		CONTROL_UNIT_OUT_PIPE: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_LD : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_MUX_CTRL : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
		CONTROL_UNIT_OUT_SUB : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		CONTROL_UNIT_OUT_SAVED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		CONTROL_UNIT_OUT_DONE : OUT STD_LOGIC);
END COMPONENT;

SIGNAL TO_STATE_REG_0,TO_STATE_REG_1,TO_STATE_REG_2,TO_STATE_REG_3,TO_STATE_REG_4,TO_STATE_REG_5,TO_STATE_REG_6,TO_STATE_REG_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_STATE_REG_0,FROM_STATE_REG_1,FROM_STATE_REG_2,FROM_STATE_REG_3,FROM_STATE_REG_4,FROM_STATE_REG_5,FROM_STATE_REG_6,FROM_STATE_REG_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_SELECTION_UNIT_0,FROM_SELECTION_UNIT_1,FROM_SELECTION_UNIT_2,FROM_SELECTION_UNIT_3,FROM_SELECTION_UNIT_4,FROM_SELECTION_UNIT_5,FROM_SELECTION_UNIT_6,FROM_SELECTION_UNIT_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_0,FROM_WINDOW_1,FROM_WINDOW_2,FROM_WINDOW_3,FROM_WINDOW_4,FROM_WINDOW_5,FROM_WINDOW_6,FROM_WINDOW_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL MASKED_INPUT_0,MASKED_INPUT_2,MASKED_INPUT_4,MASKED_INPUT_6: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_DATAPATHS_0,FROM_DATAPATHS_1,FROM_DATAPATHS_2,FROM_DATAPATHS_3,FROM_DATAPATHS_4,FROM_DATAPATHS_5,FROM_DATAPATHS_6,FROM_DATAPATHS_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_CONTROL_UNITS_0,FROM_CONTROL_UNITS_1,FROM_CONTROL_UNITS_2,FROM_CONTROL_UNITS_3,FROM_CONTROL_UNITS_4,FROM_CONTROL_UNITS_5,FROM_CONTROL_UNITS_6,FROM_CONTROL_UNITS_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL UNWINDOWED_0,UNWINDOWED_1,UNWINDOWED_2,UNWINDOWED_3,UNWINDOWED_4,UNWINDOWED_5,UNWINDOWED_6,UNWINDOWED_7: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_WINDOW_DEC_MASK : STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL UNWINDOWED_MASK, REORDERED_MASK, STATE_UPDATE_MASK : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL SELECTED_OUTPUT: STD_LOGIC_VECTOR((2*K)-1 DOWNTO 0);
SIGNAL FROM_FIRST_CU_DONE : STD_LOGIC;

BEGIN

STATE_REG_0 : n_bit_register_clear_1
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_0 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(0) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_0);
STATE_REG_1 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_1 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(1) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_1);
STATE_REG_2 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_2 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(2) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_2);
STATE_REG_3 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_3 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(3) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_3);
STATE_REG_4 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_4 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(4) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_4);
STATE_REG_5 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_5 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(5) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_5);
STATE_REG_6 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_6 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(6) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_6);
STATE_REG_7 : n_bit_register
GENERIC MAP (2*K)
PORT MAP(
												REG_IN_DATA => TO_STATE_REG_7 ,
												REG_IN_ENABLE => STATE_UPDATE_MASK(7) ,
												REG_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
												REG_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
												REG_OUT_DATA => FROM_STATE_REG_7);


MUX_SEL_UNIT_0 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_0 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_0 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_0
									);
MUX_SEL_UNIT_1 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_1 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_2 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_4 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_1
									);
MUX_SEL_UNIT_2 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_2 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_1 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_2
									);
MUX_SEL_UNIT_3 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_3 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_3 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_5 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_3
									);
MUX_SEL_UNIT_4 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_4 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_4 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_2 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_4
									);
MUX_SEL_UNIT_5 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_5 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_6 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_6 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_5
									);
MUX_SEL_UNIT_6 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_6 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_5 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_3 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_6
									);
MUX_SEL_UNIT_7 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => FROM_STATE_REG_7 ,
										MUX_3_1_IN_1 => FROM_STATE_REG_7 ,
										MUX_3_1_IN_2 => FROM_STATE_REG_7 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => FROM_SELECTION_UNIT_7
									);

MASKED_INPUT_0 <= FROM_SELECTION_UNIT_0 WHEN QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_2 <= FROM_SELECTION_UNIT_2 WHEN QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_4 <= FROM_SELECTION_UNIT_4 WHEN QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');
MASKED_INPUT_6 <= FROM_SELECTION_UNIT_6 WHEN QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF = '1' ELSE (OTHERS => '0');

FROM_WINDOW_DEC_MASK <= "1";

UNWINDOWED_MASK(0) <= QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(1) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(2) <= QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(3) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(4) <= QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(5) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(6) <= QEP_N_3_W_0_S_0_IN_MASK_FIRST_COEFF AND FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(7) <= FROM_WINDOW_DEC_MASK(0);
UNWINDOWED_MASK(7) <= FROM_WINDOW_DEC_MASK(0);
MUX_REORD_UPDATE_0 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(0 DOWNTO 0) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(0 DOWNTO 0) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(0 DOWNTO 0)
									);
MUX_REORD_UPDATE_1 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(2 DOWNTO 2) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(1 DOWNTO 1)
									);
MUX_REORD_UPDATE_2 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(2 DOWNTO 2) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(1 DOWNTO 1) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(4 DOWNTO 4) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(2 DOWNTO 2)
									);
MUX_REORD_UPDATE_3 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(3 DOWNTO 3) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(6 DOWNTO 6) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(3 DOWNTO 3)
									);
MUX_REORD_UPDATE_4 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(4 DOWNTO 4) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(1 DOWNTO 1) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(4 DOWNTO 4)
									);
MUX_REORD_UPDATE_5 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(3 DOWNTO 3) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(5 DOWNTO 5)
									);
MUX_REORD_UPDATE_6 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(6 DOWNTO 6) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(5 DOWNTO 5) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(5 DOWNTO 5) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(6 DOWNTO 6)
									);
MUX_REORD_UPDATE_7 : multiplexer_3_1 	GENERIC MAP (1)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_3_1_IN_1 => UNWINDOWED_MASK(7 DOWNTO 7) ,
										MUX_3_1_IN_2 => UNWINDOWED_MASK(7 DOWNTO 7) ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => REORDERED_MASK(7 DOWNTO 7)
									);

STATE_UPDATE_MASK(0) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(0) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(0);
STATE_UPDATE_MASK(1) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(1) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(1);
STATE_UPDATE_MASK(2) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(2) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(2);
STATE_UPDATE_MASK(3) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(3) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(3);
STATE_UPDATE_MASK(4) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(4) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(4);
STATE_UPDATE_MASK(5) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(5) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(5);
STATE_UPDATE_MASK(6) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(6) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(6);
STATE_UPDATE_MASK(7) <= QEP_N_3_W_0_S_0_IN_ENABLE_STATE_UPDATE AND FROM_FIRST_CU_DONE AND REORDERED_MASK(7) AND QEP_N_3_W_0_S_0_IN_CTRL_MASK(7);

QEP_N_3_W_0_S_0_OUT_DONE <= FROM_FIRST_CU_DONE;
CONTROL_UNIT_0 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_3_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_3_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
		CONTROL_UNIT_OUT_DONE => FROM_FIRST_CU_DONE );
CONTROL_UNIT_1 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_3_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_3_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0));
CONTROL_UNIT_2 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_3_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_3_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0));
CONTROL_UNIT_3 : control_unit PORT MAP(
		CONTROL_UNIT_IN_START =>  QEP_N_3_W_0_S_0_IN_START,
		CONTROL_UNIT_IN_OPCODE => QEP_N_3_W_0_S_0_IN_OPCODE ,
		CONTROL_UNIT_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
		CONTROL_UNIT_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
		CONTROL_UNIT_OUT_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
		CONTROL_UNIT_OUT_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
		CONTROL_UNIT_OUT_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
		CONTROL_UNIT_OUT_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
		CONTROL_UNIT_OUT_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0));

DATAPATH_0: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_0 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_1 ,
            DATAPATH_IN_SINE => QEP_N_3_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_3_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_0(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_0(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_0(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_0(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_0(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_0 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_1);
DATAPATH_1: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_2 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_3 ,
            DATAPATH_IN_SINE => QEP_N_3_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_3_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_1(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_1(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_1(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_1(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_1(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_2 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_3);
DATAPATH_2: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_4 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_5 ,
            DATAPATH_IN_SINE => QEP_N_3_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_3_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_2(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_2(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_2(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_2(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_2(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_4 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_5);
DATAPATH_3: datapath GENERIC MAP (K => K)
        PORT MAP(
            DATAPATH_IN_A => MASKED_INPUT_6 ,
            DATAPATH_IN_B => FROM_SELECTION_UNIT_7 ,
            DATAPATH_IN_SINE => QEP_N_3_W_0_S_0_IN_SIN ,
            DATAPATH_IN_COSINE => QEP_N_3_W_0_S_0_IN_COS ,
            DATAPATH_IN_PIPE => FROM_CONTROL_UNITS_3(35 DOWNTO 33) ,
            DATAPATH_IN_LD => FROM_CONTROL_UNITS_3(32 DOWNTO 30) ,
            DATAPATH_IN_MUX_CTRL => FROM_CONTROL_UNITS_3(29 DOWNTO 5) ,
            DATAPATH_IN_SUB => FROM_CONTROL_UNITS_3(4 DOWNTO 3) ,
            DATAPATH_IN_SAVED => FROM_CONTROL_UNITS_3(2 DOWNTO 0) ,
            DATAPATH_IN_CLEAR => QEP_N_3_W_0_S_0_IN_CLEAR ,
            DATAPATH_IN_CLK => QEP_N_3_W_0_S_0_IN_CLK ,
             DATAPATH_OUT_A => FROM_DATAPATHS_6 ,
            DATAPATH_OUT_B => FROM_DATAPATHS_7);

UNWINDOWED_0 <= FROM_DATAPATHS_0;
UNWINDOWED_1 <= FROM_DATAPATHS_1;
UNWINDOWED_2 <= FROM_DATAPATHS_2;
UNWINDOWED_3 <= FROM_DATAPATHS_3;
UNWINDOWED_4 <= FROM_DATAPATHS_4;
UNWINDOWED_5 <= FROM_DATAPATHS_5;
UNWINDOWED_6 <= FROM_DATAPATHS_6;
UNWINDOWED_7 <= FROM_DATAPATHS_7;

MUX_REORD_UNIT_0 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_0 ,
										MUX_3_1_IN_1 => UNWINDOWED_0 ,
										MUX_3_1_IN_2 => UNWINDOWED_0 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_0
									);
MUX_REORD_UNIT_1 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_1 ,
										MUX_3_1_IN_1 => UNWINDOWED_2 ,
										MUX_3_1_IN_2 => UNWINDOWED_2 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_1
									);
MUX_REORD_UNIT_2 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_2 ,
										MUX_3_1_IN_1 => UNWINDOWED_1 ,
										MUX_3_1_IN_2 => UNWINDOWED_4 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_2
									);
MUX_REORD_UNIT_3 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_3 ,
										MUX_3_1_IN_1 => UNWINDOWED_3 ,
										MUX_3_1_IN_2 => UNWINDOWED_6 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_3
									);
MUX_REORD_UNIT_4 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_4 ,
										MUX_3_1_IN_1 => UNWINDOWED_4 ,
										MUX_3_1_IN_2 => UNWINDOWED_1 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_4
									);
MUX_REORD_UNIT_5 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_5 ,
										MUX_3_1_IN_1 => UNWINDOWED_6 ,
										MUX_3_1_IN_2 => UNWINDOWED_3 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_5
									);
MUX_REORD_UNIT_6 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_6 ,
										MUX_3_1_IN_1 => UNWINDOWED_5 ,
										MUX_3_1_IN_2 => UNWINDOWED_5 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_6
									);
MUX_REORD_UNIT_7 : multiplexer_3_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_3_1_IN_0 => UNWINDOWED_7 ,
										MUX_3_1_IN_1 => UNWINDOWED_7 ,
										MUX_3_1_IN_2 => UNWINDOWED_7 ,
				                    			MUX_3_1_IN_SEL => QEP_N_3_W_0_S_0_IN_QTGT ,
										MUX_3_1_OUT_RES => TO_STATE_REG_7
									);

MUX_OUTPUT_SELECTION : multiplexer_8_1 	GENERIC MAP (2*K)
									PORT MAP (
										MUX_8_1_IN_0 => FROM_STATE_REG_0 ,
										MUX_8_1_IN_1 => FROM_STATE_REG_1 ,
										MUX_8_1_IN_2 => FROM_STATE_REG_2 ,
										MUX_8_1_IN_3 => FROM_STATE_REG_3 ,
										MUX_8_1_IN_4 => FROM_STATE_REG_4 ,
										MUX_8_1_IN_5 => FROM_STATE_REG_5 ,
										MUX_8_1_IN_6 => FROM_STATE_REG_6 ,
										MUX_8_1_IN_7 => FROM_STATE_REG_7 ,
				                    			MUX_8_1_IN_SEL => QEP_N_3_W_0_S_0_IN_OUT_STATE_SEL ,
										MUX_8_1_OUT_RES => SELECTED_OUTPUT
									);
MUX_REAL_IMAG_SELECTION : multiplexer_2_1 GENERIC MAP (K => K)
									PORT MAP (
										MUX_2_1_IN_0 => SELECTED_OUTPUT((2*K-1) DOWNTO K),
										MUX_2_1_IN_1 => SELECTED_OUTPUT((K-1) DOWNTO 0),
				                    			MUX_2_1_IN_SEL => QEP_N_3_W_0_S_0_IN_REAL_IMAG_SEL ,
										MUX_2_1_OUT_RES => QEP_N_3_W_0_S_0_OUT_DATA
									);

END generated;