library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_2_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_2_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_2_1_IN_SEL : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		MUX_2_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_2_1 IS

BEGIN

	MUX_2_1_OUT_RES <= 
				MUX_2_1_IN_0 WHEN MUX_2_1_IN_SEL = "0" ELSE
				MUX_2_1_IN_1 WHEN MUX_2_1_IN_SEL = "1" ELSE
				(OTHERS => '0');


END behavioral;