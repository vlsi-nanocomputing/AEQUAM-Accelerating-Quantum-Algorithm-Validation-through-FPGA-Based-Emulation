library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_9_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_9_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_9_1_IN_SEL : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		MUX_9_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_9_1 IS

BEGIN

	MUX_9_1_OUT_RES <= 
				MUX_9_1_IN_0 WHEN MUX_9_1_IN_SEL = "0000" ELSE
				MUX_9_1_IN_1 WHEN MUX_9_1_IN_SEL = "0001" ELSE
				MUX_9_1_IN_2 WHEN MUX_9_1_IN_SEL = "0010" ELSE
				MUX_9_1_IN_3 WHEN MUX_9_1_IN_SEL = "0011" ELSE
				MUX_9_1_IN_4 WHEN MUX_9_1_IN_SEL = "0100" ELSE
				MUX_9_1_IN_5 WHEN MUX_9_1_IN_SEL = "0101" ELSE
				MUX_9_1_IN_6 WHEN MUX_9_1_IN_SEL = "0110" ELSE
				MUX_9_1_IN_7 WHEN MUX_9_1_IN_SEL = "0111" ELSE
				MUX_9_1_IN_8 WHEN MUX_9_1_IN_SEL = "1000" ELSE
				(OTHERS => '0');


END behavioral;