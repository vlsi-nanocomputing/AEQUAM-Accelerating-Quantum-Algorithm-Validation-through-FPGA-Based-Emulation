library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
ENTITY multiplexer_32_1 IS 
	GENERIC (K : INTEGER := 20);
	PORT (
		MUX_32_1_IN_0 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_1 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_2 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_3 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_4 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_5 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_6 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_7 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_8 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_9 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_10 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_11 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_12 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_13 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_14 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_15 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_16 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_17 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_18 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_19 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_20 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_21 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_22 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_23 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_24 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_25 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_26 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_27 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_28 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_29 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_30 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_31 : IN STD_LOGIC_VECTOR (K-1 DOWNTO 0);
		MUX_32_1_IN_SEL : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		MUX_32_1_OUT_RES : OUT STD_LOGIC_VECTOR (K-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE behavioral OF multiplexer_32_1 IS

BEGIN

	MUX_32_1_OUT_RES <= 
				MUX_32_1_IN_0 WHEN MUX_32_1_IN_SEL = "00000" ELSE
				MUX_32_1_IN_1 WHEN MUX_32_1_IN_SEL = "00001" ELSE
				MUX_32_1_IN_2 WHEN MUX_32_1_IN_SEL = "00010" ELSE
				MUX_32_1_IN_3 WHEN MUX_32_1_IN_SEL = "00011" ELSE
				MUX_32_1_IN_4 WHEN MUX_32_1_IN_SEL = "00100" ELSE
				MUX_32_1_IN_5 WHEN MUX_32_1_IN_SEL = "00101" ELSE
				MUX_32_1_IN_6 WHEN MUX_32_1_IN_SEL = "00110" ELSE
				MUX_32_1_IN_7 WHEN MUX_32_1_IN_SEL = "00111" ELSE
				MUX_32_1_IN_8 WHEN MUX_32_1_IN_SEL = "01000" ELSE
				MUX_32_1_IN_9 WHEN MUX_32_1_IN_SEL = "01001" ELSE
				MUX_32_1_IN_10 WHEN MUX_32_1_IN_SEL = "01010" ELSE
				MUX_32_1_IN_11 WHEN MUX_32_1_IN_SEL = "01011" ELSE
				MUX_32_1_IN_12 WHEN MUX_32_1_IN_SEL = "01100" ELSE
				MUX_32_1_IN_13 WHEN MUX_32_1_IN_SEL = "01101" ELSE
				MUX_32_1_IN_14 WHEN MUX_32_1_IN_SEL = "01110" ELSE
				MUX_32_1_IN_15 WHEN MUX_32_1_IN_SEL = "01111" ELSE
				MUX_32_1_IN_16 WHEN MUX_32_1_IN_SEL = "10000" ELSE
				MUX_32_1_IN_17 WHEN MUX_32_1_IN_SEL = "10001" ELSE
				MUX_32_1_IN_18 WHEN MUX_32_1_IN_SEL = "10010" ELSE
				MUX_32_1_IN_19 WHEN MUX_32_1_IN_SEL = "10011" ELSE
				MUX_32_1_IN_20 WHEN MUX_32_1_IN_SEL = "10100" ELSE
				MUX_32_1_IN_21 WHEN MUX_32_1_IN_SEL = "10101" ELSE
				MUX_32_1_IN_22 WHEN MUX_32_1_IN_SEL = "10110" ELSE
				MUX_32_1_IN_23 WHEN MUX_32_1_IN_SEL = "10111" ELSE
				MUX_32_1_IN_24 WHEN MUX_32_1_IN_SEL = "11000" ELSE
				MUX_32_1_IN_25 WHEN MUX_32_1_IN_SEL = "11001" ELSE
				MUX_32_1_IN_26 WHEN MUX_32_1_IN_SEL = "11010" ELSE
				MUX_32_1_IN_27 WHEN MUX_32_1_IN_SEL = "11011" ELSE
				MUX_32_1_IN_28 WHEN MUX_32_1_IN_SEL = "11100" ELSE
				MUX_32_1_IN_29 WHEN MUX_32_1_IN_SEL = "11101" ELSE
				MUX_32_1_IN_30 WHEN MUX_32_1_IN_SEL = "11110" ELSE
				MUX_32_1_IN_31 WHEN MUX_32_1_IN_SEL = "11111" ELSE
				(OTHERS => '0');


END behavioral;